module  M_TWIDLE_8_bit #(parameter SIZE =10, word_length_tw = 8) (
    input            clk,
    input            en_rd, 
    input   [10:0]   rd_ptr_angle,
    input            en_modf, 

    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );


reg signed [word_length_tw-1:0]  cos  [511:0];
reg signed [word_length_tw-1:0]  sin  [511:0];

reg signed [word_length_tw-1:0]  m_cos  [511:0];
reg signed [word_length_tw-1:0]  m_sin  [511:0];

reg signed [word_length_tw-1:0]  cos_temp;
reg signed [word_length_tw-1:0]  sin_temp;

reg signed [word_length_tw-1:0]  m_cos_temp;
reg signed [word_length_tw-1:0]  m_sin_temp;


//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & ~ en_modf ) begin
                  cos_temp           <= cos   [rd_ptr_angle];
                  sin_temp           <= sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & en_modf ) begin
                  m_cos_temp           <= m_cos   [rd_ptr_angle];
                  m_sin_temp           <= m_sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(*) begin 
             if (en_modf ) begin
                  cos_data           <= m_cos_temp;
                  sin_data           <= m_sin_temp;
             end else begin
                  cos_data           <= cos_temp;
                  sin_data           <= sin_temp;
             end
        end
//----------------------------------------------------------------------------------------
initial begin
   sin[0]  =  8'b00000000;     //0pi/512
   cos[0]  =  8'b01000000;     //0pi/512
   sin[1]  =  8'b00000000;     //1pi/512
   cos[1]  =  8'b00111111;     //1pi/512
   sin[2]  =  8'b11111111;     //2pi/512
   cos[2]  =  8'b00111111;     //2pi/512
   sin[3]  =  8'b11111111;     //3pi/512
   cos[3]  =  8'b00111111;     //3pi/512
   sin[4]  =  8'b11111110;     //4pi/512
   cos[4]  =  8'b00111111;     //4pi/512
   sin[5]  =  8'b11111110;     //5pi/512
   cos[5]  =  8'b00111111;     //5pi/512
   sin[6]  =  8'b11111110;     //6pi/512
   cos[6]  =  8'b00111111;     //6pi/512
   sin[7]  =  8'b11111101;     //7pi/512
   cos[7]  =  8'b00111111;     //7pi/512
   sin[8]  =  8'b11111101;     //8pi/512
   cos[8]  =  8'b00111111;     //8pi/512
   sin[9]  =  8'b11111100;     //9pi/512
   cos[9]  =  8'b00111111;     //9pi/512
   sin[10]  =  8'b11111100;     //10pi/512
   cos[10]  =  8'b00111111;     //10pi/512
   sin[11]  =  8'b11111100;     //11pi/512
   cos[11]  =  8'b00111111;     //11pi/512
   sin[12]  =  8'b11111011;     //12pi/512
   cos[12]  =  8'b00111111;     //12pi/512
   sin[13]  =  8'b11111011;     //13pi/512
   cos[13]  =  8'b00111111;     //13pi/512
   sin[14]  =  8'b11111011;     //14pi/512
   cos[14]  =  8'b00111111;     //14pi/512
   sin[15]  =  8'b11111010;     //15pi/512
   cos[15]  =  8'b00111111;     //15pi/512
   sin[16]  =  8'b11111010;     //16pi/512
   cos[16]  =  8'b00111111;     //16pi/512
   sin[17]  =  8'b11111001;     //17pi/512
   cos[17]  =  8'b00111111;     //17pi/512
   sin[18]  =  8'b11111001;     //18pi/512
   cos[18]  =  8'b00111111;     //18pi/512
   sin[19]  =  8'b11111001;     //19pi/512
   cos[19]  =  8'b00111111;     //19pi/512
   sin[20]  =  8'b11111000;     //20pi/512
   cos[20]  =  8'b00111111;     //20pi/512
   sin[21]  =  8'b11111000;     //21pi/512
   cos[21]  =  8'b00111111;     //21pi/512
   sin[22]  =  8'b11110111;     //22pi/512
   cos[22]  =  8'b00111111;     //22pi/512
   sin[23]  =  8'b11110111;     //23pi/512
   cos[23]  =  8'b00111111;     //23pi/512
   sin[24]  =  8'b11110111;     //24pi/512
   cos[24]  =  8'b00111111;     //24pi/512
   sin[25]  =  8'b11110110;     //25pi/512
   cos[25]  =  8'b00111111;     //25pi/512
   sin[26]  =  8'b11110110;     //26pi/512
   cos[26]  =  8'b00111111;     //26pi/512
   sin[27]  =  8'b11110101;     //27pi/512
   cos[27]  =  8'b00111111;     //27pi/512
   sin[28]  =  8'b11110101;     //28pi/512
   cos[28]  =  8'b00111111;     //28pi/512
   sin[29]  =  8'b11110101;     //29pi/512
   cos[29]  =  8'b00111110;     //29pi/512
   sin[30]  =  8'b11110100;     //30pi/512
   cos[30]  =  8'b00111110;     //30pi/512
   sin[31]  =  8'b11110100;     //31pi/512
   cos[31]  =  8'b00111110;     //31pi/512
   sin[32]  =  8'b11110100;     //32pi/512
   cos[32]  =  8'b00111110;     //32pi/512
   sin[33]  =  8'b11110011;     //33pi/512
   cos[33]  =  8'b00111110;     //33pi/512
   sin[34]  =  8'b11110011;     //34pi/512
   cos[34]  =  8'b00111110;     //34pi/512
   sin[35]  =  8'b11110010;     //35pi/512
   cos[35]  =  8'b00111110;     //35pi/512
   sin[36]  =  8'b11110010;     //36pi/512
   cos[36]  =  8'b00111110;     //36pi/512
   sin[37]  =  8'b11110010;     //37pi/512
   cos[37]  =  8'b00111110;     //37pi/512
   sin[38]  =  8'b11110001;     //38pi/512
   cos[38]  =  8'b00111110;     //38pi/512
   sin[39]  =  8'b11110001;     //39pi/512
   cos[39]  =  8'b00111110;     //39pi/512
   sin[40]  =  8'b11110000;     //40pi/512
   cos[40]  =  8'b00111110;     //40pi/512
   sin[41]  =  8'b11110000;     //41pi/512
   cos[41]  =  8'b00111101;     //41pi/512
   sin[42]  =  8'b11110000;     //42pi/512
   cos[42]  =  8'b00111101;     //42pi/512
   sin[43]  =  8'b11101111;     //43pi/512
   cos[43]  =  8'b00111101;     //43pi/512
   sin[44]  =  8'b11101111;     //44pi/512
   cos[44]  =  8'b00111101;     //44pi/512
   sin[45]  =  8'b11101111;     //45pi/512
   cos[45]  =  8'b00111101;     //45pi/512
   sin[46]  =  8'b11101110;     //46pi/512
   cos[46]  =  8'b00111101;     //46pi/512
   sin[47]  =  8'b11101110;     //47pi/512
   cos[47]  =  8'b00111101;     //47pi/512
   sin[48]  =  8'b11101101;     //48pi/512
   cos[48]  =  8'b00111101;     //48pi/512
   sin[49]  =  8'b11101101;     //49pi/512
   cos[49]  =  8'b00111101;     //49pi/512
   sin[50]  =  8'b11101101;     //50pi/512
   cos[50]  =  8'b00111101;     //50pi/512
   sin[51]  =  8'b11101100;     //51pi/512
   cos[51]  =  8'b00111100;     //51pi/512
   sin[52]  =  8'b11101100;     //52pi/512
   cos[52]  =  8'b00111100;     //52pi/512
   sin[53]  =  8'b11101100;     //53pi/512
   cos[53]  =  8'b00111100;     //53pi/512
   sin[54]  =  8'b11101011;     //54pi/512
   cos[54]  =  8'b00111100;     //54pi/512
   sin[55]  =  8'b11101011;     //55pi/512
   cos[55]  =  8'b00111100;     //55pi/512
   sin[56]  =  8'b11101010;     //56pi/512
   cos[56]  =  8'b00111100;     //56pi/512
   sin[57]  =  8'b11101010;     //57pi/512
   cos[57]  =  8'b00111100;     //57pi/512
   sin[58]  =  8'b11101010;     //58pi/512
   cos[58]  =  8'b00111011;     //58pi/512
   sin[59]  =  8'b11101001;     //59pi/512
   cos[59]  =  8'b00111011;     //59pi/512
   sin[60]  =  8'b11101001;     //60pi/512
   cos[60]  =  8'b00111011;     //60pi/512
   sin[61]  =  8'b11101001;     //61pi/512
   cos[61]  =  8'b00111011;     //61pi/512
   sin[62]  =  8'b11101000;     //62pi/512
   cos[62]  =  8'b00111011;     //62pi/512
   sin[63]  =  8'b11101000;     //63pi/512
   cos[63]  =  8'b00111011;     //63pi/512
   sin[64]  =  8'b11101000;     //64pi/512
   cos[64]  =  8'b00111011;     //64pi/512
   sin[65]  =  8'b11100111;     //65pi/512
   cos[65]  =  8'b00111010;     //65pi/512
   sin[66]  =  8'b11100111;     //66pi/512
   cos[66]  =  8'b00111010;     //66pi/512
   sin[67]  =  8'b11100110;     //67pi/512
   cos[67]  =  8'b00111010;     //67pi/512
   sin[68]  =  8'b11100110;     //68pi/512
   cos[68]  =  8'b00111010;     //68pi/512
   sin[69]  =  8'b11100110;     //69pi/512
   cos[69]  =  8'b00111010;     //69pi/512
   sin[70]  =  8'b11100101;     //70pi/512
   cos[70]  =  8'b00111010;     //70pi/512
   sin[71]  =  8'b11100101;     //71pi/512
   cos[71]  =  8'b00111010;     //71pi/512
   sin[72]  =  8'b11100101;     //72pi/512
   cos[72]  =  8'b00111001;     //72pi/512
   sin[73]  =  8'b11100100;     //73pi/512
   cos[73]  =  8'b00111001;     //73pi/512
   sin[74]  =  8'b11100100;     //74pi/512
   cos[74]  =  8'b00111001;     //74pi/512
   sin[75]  =  8'b11100100;     //75pi/512
   cos[75]  =  8'b00111001;     //75pi/512
   sin[76]  =  8'b11100011;     //76pi/512
   cos[76]  =  8'b00111001;     //76pi/512
   sin[77]  =  8'b11100011;     //77pi/512
   cos[77]  =  8'b00111000;     //77pi/512
   sin[78]  =  8'b11100011;     //78pi/512
   cos[78]  =  8'b00111000;     //78pi/512
   sin[79]  =  8'b11100010;     //79pi/512
   cos[79]  =  8'b00111000;     //79pi/512
   sin[80]  =  8'b11100010;     //80pi/512
   cos[80]  =  8'b00111000;     //80pi/512
   sin[81]  =  8'b11100001;     //81pi/512
   cos[81]  =  8'b00111000;     //81pi/512
   sin[82]  =  8'b11100001;     //82pi/512
   cos[82]  =  8'b00111000;     //82pi/512
   sin[83]  =  8'b11100001;     //83pi/512
   cos[83]  =  8'b00110111;     //83pi/512
   sin[84]  =  8'b11100000;     //84pi/512
   cos[84]  =  8'b00110111;     //84pi/512
   sin[85]  =  8'b11100000;     //85pi/512
   cos[85]  =  8'b00110111;     //85pi/512
   sin[86]  =  8'b11100000;     //86pi/512
   cos[86]  =  8'b00110111;     //86pi/512
   sin[87]  =  8'b11011111;     //87pi/512
   cos[87]  =  8'b00110111;     //87pi/512
   sin[88]  =  8'b11011111;     //88pi/512
   cos[88]  =  8'b00110110;     //88pi/512
   sin[89]  =  8'b11011111;     //89pi/512
   cos[89]  =  8'b00110110;     //89pi/512
   sin[90]  =  8'b11011110;     //90pi/512
   cos[90]  =  8'b00110110;     //90pi/512
   sin[91]  =  8'b11011110;     //91pi/512
   cos[91]  =  8'b00110110;     //91pi/512
   sin[92]  =  8'b11011110;     //92pi/512
   cos[92]  =  8'b00110110;     //92pi/512
   sin[93]  =  8'b11011101;     //93pi/512
   cos[93]  =  8'b00110101;     //93pi/512
   sin[94]  =  8'b11011101;     //94pi/512
   cos[94]  =  8'b00110101;     //94pi/512
   sin[95]  =  8'b11011101;     //95pi/512
   cos[95]  =  8'b00110101;     //95pi/512
   sin[96]  =  8'b11011100;     //96pi/512
   cos[96]  =  8'b00110101;     //96pi/512
   sin[97]  =  8'b11011100;     //97pi/512
   cos[97]  =  8'b00110100;     //97pi/512
   sin[98]  =  8'b11011100;     //98pi/512
   cos[98]  =  8'b00110100;     //98pi/512
   sin[99]  =  8'b11011011;     //99pi/512
   cos[99]  =  8'b00110100;     //99pi/512
   sin[100]  =  8'b11011011;     //100pi/512
   cos[100]  =  8'b00110100;     //100pi/512
   sin[101]  =  8'b11011011;     //101pi/512
   cos[101]  =  8'b00110100;     //101pi/512
   sin[102]  =  8'b11011011;     //102pi/512
   cos[102]  =  8'b00110011;     //102pi/512
   sin[103]  =  8'b11011010;     //103pi/512
   cos[103]  =  8'b00110011;     //103pi/512
   sin[104]  =  8'b11011010;     //104pi/512
   cos[104]  =  8'b00110011;     //104pi/512
   sin[105]  =  8'b11011010;     //105pi/512
   cos[105]  =  8'b00110011;     //105pi/512
   sin[106]  =  8'b11011001;     //106pi/512
   cos[106]  =  8'b00110010;     //106pi/512
   sin[107]  =  8'b11011001;     //107pi/512
   cos[107]  =  8'b00110010;     //107pi/512
   sin[108]  =  8'b11011001;     //108pi/512
   cos[108]  =  8'b00110010;     //108pi/512
   sin[109]  =  8'b11011000;     //109pi/512
   cos[109]  =  8'b00110010;     //109pi/512
   sin[110]  =  8'b11011000;     //110pi/512
   cos[110]  =  8'b00110001;     //110pi/512
   sin[111]  =  8'b11011000;     //111pi/512
   cos[111]  =  8'b00110001;     //111pi/512
   sin[112]  =  8'b11010111;     //112pi/512
   cos[112]  =  8'b00110001;     //112pi/512
   sin[113]  =  8'b11010111;     //113pi/512
   cos[113]  =  8'b00110001;     //113pi/512
   sin[114]  =  8'b11010111;     //114pi/512
   cos[114]  =  8'b00110000;     //114pi/512
   sin[115]  =  8'b11010110;     //115pi/512
   cos[115]  =  8'b00110000;     //115pi/512
   sin[116]  =  8'b11010110;     //116pi/512
   cos[116]  =  8'b00110000;     //116pi/512
   sin[117]  =  8'b11010110;     //117pi/512
   cos[117]  =  8'b00110000;     //117pi/512
   sin[118]  =  8'b11010110;     //118pi/512
   cos[118]  =  8'b00101111;     //118pi/512
   sin[119]  =  8'b11010101;     //119pi/512
   cos[119]  =  8'b00101111;     //119pi/512
   sin[120]  =  8'b11010101;     //120pi/512
   cos[120]  =  8'b00101111;     //120pi/512
   sin[121]  =  8'b11010101;     //121pi/512
   cos[121]  =  8'b00101111;     //121pi/512
   sin[122]  =  8'b11010100;     //122pi/512
   cos[122]  =  8'b00101110;     //122pi/512
   sin[123]  =  8'b11010100;     //123pi/512
   cos[123]  =  8'b00101110;     //123pi/512
   sin[124]  =  8'b11010100;     //124pi/512
   cos[124]  =  8'b00101110;     //124pi/512
   sin[125]  =  8'b11010100;     //125pi/512
   cos[125]  =  8'b00101110;     //125pi/512
   sin[126]  =  8'b11010011;     //126pi/512
   cos[126]  =  8'b00101101;     //126pi/512
   sin[127]  =  8'b11010011;     //127pi/512
   cos[127]  =  8'b00101101;     //127pi/512
   sin[128]  =  8'b11010011;     //128pi/512
   cos[128]  =  8'b00101101;     //128pi/512
   sin[129]  =  8'b11010010;     //129pi/512
   cos[129]  =  8'b00101100;     //129pi/512
   sin[130]  =  8'b11010010;     //130pi/512
   cos[130]  =  8'b00101100;     //130pi/512
   sin[131]  =  8'b11010010;     //131pi/512
   cos[131]  =  8'b00101100;     //131pi/512
   sin[132]  =  8'b11010010;     //132pi/512
   cos[132]  =  8'b00101100;     //132pi/512
   sin[133]  =  8'b11010001;     //133pi/512
   cos[133]  =  8'b00101011;     //133pi/512
   sin[134]  =  8'b11010001;     //134pi/512
   cos[134]  =  8'b00101011;     //134pi/512
   sin[135]  =  8'b11010001;     //135pi/512
   cos[135]  =  8'b00101011;     //135pi/512
   sin[136]  =  8'b11010001;     //136pi/512
   cos[136]  =  8'b00101010;     //136pi/512
   sin[137]  =  8'b11010000;     //137pi/512
   cos[137]  =  8'b00101010;     //137pi/512
   sin[138]  =  8'b11010000;     //138pi/512
   cos[138]  =  8'b00101010;     //138pi/512
   sin[139]  =  8'b11010000;     //139pi/512
   cos[139]  =  8'b00101010;     //139pi/512
   sin[140]  =  8'b11010000;     //140pi/512
   cos[140]  =  8'b00101001;     //140pi/512
   sin[141]  =  8'b11001111;     //141pi/512
   cos[141]  =  8'b00101001;     //141pi/512
   sin[142]  =  8'b11001111;     //142pi/512
   cos[142]  =  8'b00101001;     //142pi/512
   sin[143]  =  8'b11001111;     //143pi/512
   cos[143]  =  8'b00101000;     //143pi/512
   sin[144]  =  8'b11001111;     //144pi/512
   cos[144]  =  8'b00101000;     //144pi/512
   sin[145]  =  8'b11001110;     //145pi/512
   cos[145]  =  8'b00101000;     //145pi/512
   sin[146]  =  8'b11001110;     //146pi/512
   cos[146]  =  8'b00100111;     //146pi/512
   sin[147]  =  8'b11001110;     //147pi/512
   cos[147]  =  8'b00100111;     //147pi/512
   sin[148]  =  8'b11001110;     //148pi/512
   cos[148]  =  8'b00100111;     //148pi/512
   sin[149]  =  8'b11001101;     //149pi/512
   cos[149]  =  8'b00100111;     //149pi/512
   sin[150]  =  8'b11001101;     //150pi/512
   cos[150]  =  8'b00100110;     //150pi/512
   sin[151]  =  8'b11001101;     //151pi/512
   cos[151]  =  8'b00100110;     //151pi/512
   sin[152]  =  8'b11001101;     //152pi/512
   cos[152]  =  8'b00100110;     //152pi/512
   sin[153]  =  8'b11001100;     //153pi/512
   cos[153]  =  8'b00100101;     //153pi/512
   sin[154]  =  8'b11001100;     //154pi/512
   cos[154]  =  8'b00100101;     //154pi/512
   sin[155]  =  8'b11001100;     //155pi/512
   cos[155]  =  8'b00100101;     //155pi/512
   sin[156]  =  8'b11001100;     //156pi/512
   cos[156]  =  8'b00100100;     //156pi/512
   sin[157]  =  8'b11001011;     //157pi/512
   cos[157]  =  8'b00100100;     //157pi/512
   sin[158]  =  8'b11001011;     //158pi/512
   cos[158]  =  8'b00100100;     //158pi/512
   sin[159]  =  8'b11001011;     //159pi/512
   cos[159]  =  8'b00100011;     //159pi/512
   sin[160]  =  8'b11001011;     //160pi/512
   cos[160]  =  8'b00100011;     //160pi/512
   sin[161]  =  8'b11001011;     //161pi/512
   cos[161]  =  8'b00100011;     //161pi/512
   sin[162]  =  8'b11001010;     //162pi/512
   cos[162]  =  8'b00100010;     //162pi/512
   sin[163]  =  8'b11001010;     //163pi/512
   cos[163]  =  8'b00100010;     //163pi/512
   sin[164]  =  8'b11001010;     //164pi/512
   cos[164]  =  8'b00100010;     //164pi/512
   sin[165]  =  8'b11001010;     //165pi/512
   cos[165]  =  8'b00100001;     //165pi/512
   sin[166]  =  8'b11001010;     //166pi/512
   cos[166]  =  8'b00100001;     //166pi/512
   sin[167]  =  8'b11001001;     //167pi/512
   cos[167]  =  8'b00100001;     //167pi/512
   sin[168]  =  8'b11001001;     //168pi/512
   cos[168]  =  8'b00100000;     //168pi/512
   sin[169]  =  8'b11001001;     //169pi/512
   cos[169]  =  8'b00100000;     //169pi/512
   sin[170]  =  8'b11001001;     //170pi/512
   cos[170]  =  8'b00100000;     //170pi/512
   sin[171]  =  8'b11001001;     //171pi/512
   cos[171]  =  8'b00011111;     //171pi/512
   sin[172]  =  8'b11001000;     //172pi/512
   cos[172]  =  8'b00011111;     //172pi/512
   sin[173]  =  8'b11001000;     //173pi/512
   cos[173]  =  8'b00011111;     //173pi/512
   sin[174]  =  8'b11001000;     //174pi/512
   cos[174]  =  8'b00011110;     //174pi/512
   sin[175]  =  8'b11001000;     //175pi/512
   cos[175]  =  8'b00011110;     //175pi/512
   sin[176]  =  8'b11001000;     //176pi/512
   cos[176]  =  8'b00011110;     //176pi/512
   sin[177]  =  8'b11000111;     //177pi/512
   cos[177]  =  8'b00011101;     //177pi/512
   sin[178]  =  8'b11000111;     //178pi/512
   cos[178]  =  8'b00011101;     //178pi/512
   sin[179]  =  8'b11000111;     //179pi/512
   cos[179]  =  8'b00011101;     //179pi/512
   sin[180]  =  8'b11000111;     //180pi/512
   cos[180]  =  8'b00011100;     //180pi/512
   sin[181]  =  8'b11000111;     //181pi/512
   cos[181]  =  8'b00011100;     //181pi/512
   sin[182]  =  8'b11000110;     //182pi/512
   cos[182]  =  8'b00011100;     //182pi/512
   sin[183]  =  8'b11000110;     //183pi/512
   cos[183]  =  8'b00011011;     //183pi/512
   sin[184]  =  8'b11000110;     //184pi/512
   cos[184]  =  8'b00011011;     //184pi/512
   sin[185]  =  8'b11000110;     //185pi/512
   cos[185]  =  8'b00011011;     //185pi/512
   sin[186]  =  8'b11000110;     //186pi/512
   cos[186]  =  8'b00011010;     //186pi/512
   sin[187]  =  8'b11000110;     //187pi/512
   cos[187]  =  8'b00011010;     //187pi/512
   sin[188]  =  8'b11000101;     //188pi/512
   cos[188]  =  8'b00011001;     //188pi/512
   sin[189]  =  8'b11000101;     //189pi/512
   cos[189]  =  8'b00011001;     //189pi/512
   sin[190]  =  8'b11000101;     //190pi/512
   cos[190]  =  8'b00011001;     //190pi/512
   sin[191]  =  8'b11000101;     //191pi/512
   cos[191]  =  8'b00011000;     //191pi/512
   sin[192]  =  8'b11000101;     //192pi/512
   cos[192]  =  8'b00011000;     //192pi/512
   sin[193]  =  8'b11000101;     //193pi/512
   cos[193]  =  8'b00011000;     //193pi/512
   sin[194]  =  8'b11000101;     //194pi/512
   cos[194]  =  8'b00010111;     //194pi/512
   sin[195]  =  8'b11000100;     //195pi/512
   cos[195]  =  8'b00010111;     //195pi/512
   sin[196]  =  8'b11000100;     //196pi/512
   cos[196]  =  8'b00010111;     //196pi/512
   sin[197]  =  8'b11000100;     //197pi/512
   cos[197]  =  8'b00010110;     //197pi/512
   sin[198]  =  8'b11000100;     //198pi/512
   cos[198]  =  8'b00010110;     //198pi/512
   sin[199]  =  8'b11000100;     //199pi/512
   cos[199]  =  8'b00010101;     //199pi/512
   sin[200]  =  8'b11000100;     //200pi/512
   cos[200]  =  8'b00010101;     //200pi/512
   sin[201]  =  8'b11000100;     //201pi/512
   cos[201]  =  8'b00010101;     //201pi/512
   sin[202]  =  8'b11000011;     //202pi/512
   cos[202]  =  8'b00010100;     //202pi/512
   sin[203]  =  8'b11000011;     //203pi/512
   cos[203]  =  8'b00010100;     //203pi/512
   sin[204]  =  8'b11000011;     //204pi/512
   cos[204]  =  8'b00010100;     //204pi/512
   sin[205]  =  8'b11000011;     //205pi/512
   cos[205]  =  8'b00010011;     //205pi/512
   sin[206]  =  8'b11000011;     //206pi/512
   cos[206]  =  8'b00010011;     //206pi/512
   sin[207]  =  8'b11000011;     //207pi/512
   cos[207]  =  8'b00010010;     //207pi/512
   sin[208]  =  8'b11000011;     //208pi/512
   cos[208]  =  8'b00010010;     //208pi/512
   sin[209]  =  8'b11000011;     //209pi/512
   cos[209]  =  8'b00010010;     //209pi/512
   sin[210]  =  8'b11000011;     //210pi/512
   cos[210]  =  8'b00010001;     //210pi/512
   sin[211]  =  8'b11000010;     //211pi/512
   cos[211]  =  8'b00010001;     //211pi/512
   sin[212]  =  8'b11000010;     //212pi/512
   cos[212]  =  8'b00010001;     //212pi/512
   sin[213]  =  8'b11000010;     //213pi/512
   cos[213]  =  8'b00010000;     //213pi/512
   sin[214]  =  8'b11000010;     //214pi/512
   cos[214]  =  8'b00010000;     //214pi/512
   sin[215]  =  8'b11000010;     //215pi/512
   cos[215]  =  8'b00001111;     //215pi/512
   sin[216]  =  8'b11000010;     //216pi/512
   cos[216]  =  8'b00001111;     //216pi/512
   sin[217]  =  8'b11000010;     //217pi/512
   cos[217]  =  8'b00001111;     //217pi/512
   sin[218]  =  8'b11000010;     //218pi/512
   cos[218]  =  8'b00001110;     //218pi/512
   sin[219]  =  8'b11000010;     //219pi/512
   cos[219]  =  8'b00001110;     //219pi/512
   sin[220]  =  8'b11000010;     //220pi/512
   cos[220]  =  8'b00001110;     //220pi/512
   sin[221]  =  8'b11000001;     //221pi/512
   cos[221]  =  8'b00001101;     //221pi/512
   sin[222]  =  8'b11000001;     //222pi/512
   cos[222]  =  8'b00001101;     //222pi/512
   sin[223]  =  8'b11000001;     //223pi/512
   cos[223]  =  8'b00001100;     //223pi/512
   sin[224]  =  8'b11000001;     //224pi/512
   cos[224]  =  8'b00001100;     //224pi/512
   sin[225]  =  8'b11000001;     //225pi/512
   cos[225]  =  8'b00001100;     //225pi/512
   sin[226]  =  8'b11000001;     //226pi/512
   cos[226]  =  8'b00001011;     //226pi/512
   sin[227]  =  8'b11000001;     //227pi/512
   cos[227]  =  8'b00001011;     //227pi/512
   sin[228]  =  8'b11000001;     //228pi/512
   cos[228]  =  8'b00001010;     //228pi/512
   sin[229]  =  8'b11000001;     //229pi/512
   cos[229]  =  8'b00001010;     //229pi/512
   sin[230]  =  8'b11000001;     //230pi/512
   cos[230]  =  8'b00001010;     //230pi/512
   sin[231]  =  8'b11000001;     //231pi/512
   cos[231]  =  8'b00001001;     //231pi/512
   sin[232]  =  8'b11000001;     //232pi/512
   cos[232]  =  8'b00001001;     //232pi/512
   sin[233]  =  8'b11000001;     //233pi/512
   cos[233]  =  8'b00001001;     //233pi/512
   sin[234]  =  8'b11000001;     //234pi/512
   cos[234]  =  8'b00001000;     //234pi/512
   sin[235]  =  8'b11000001;     //235pi/512
   cos[235]  =  8'b00001000;     //235pi/512
   sin[236]  =  8'b11000000;     //236pi/512
   cos[236]  =  8'b00000111;     //236pi/512
   sin[237]  =  8'b11000000;     //237pi/512
   cos[237]  =  8'b00000111;     //237pi/512
   sin[238]  =  8'b11000000;     //238pi/512
   cos[238]  =  8'b00000111;     //238pi/512
   sin[239]  =  8'b11000000;     //239pi/512
   cos[239]  =  8'b00000110;     //239pi/512
   sin[240]  =  8'b11000000;     //240pi/512
   cos[240]  =  8'b00000110;     //240pi/512
   sin[241]  =  8'b11000000;     //241pi/512
   cos[241]  =  8'b00000101;     //241pi/512
   sin[242]  =  8'b11000000;     //242pi/512
   cos[242]  =  8'b00000101;     //242pi/512
   sin[243]  =  8'b11000000;     //243pi/512
   cos[243]  =  8'b00000101;     //243pi/512
   sin[244]  =  8'b11000000;     //244pi/512
   cos[244]  =  8'b00000100;     //244pi/512
   sin[245]  =  8'b11000000;     //245pi/512
   cos[245]  =  8'b00000100;     //245pi/512
   sin[246]  =  8'b11000000;     //246pi/512
   cos[246]  =  8'b00000011;     //246pi/512
   sin[247]  =  8'b11000000;     //247pi/512
   cos[247]  =  8'b00000011;     //247pi/512
   sin[248]  =  8'b11000000;     //248pi/512
   cos[248]  =  8'b00000011;     //248pi/512
   sin[249]  =  8'b11000000;     //249pi/512
   cos[249]  =  8'b00000010;     //249pi/512
   sin[250]  =  8'b11000000;     //250pi/512
   cos[250]  =  8'b00000010;     //250pi/512
   sin[251]  =  8'b11000000;     //251pi/512
   cos[251]  =  8'b00000001;     //251pi/512
   sin[252]  =  8'b11000000;     //252pi/512
   cos[252]  =  8'b00000001;     //252pi/512
   sin[253]  =  8'b11000000;     //253pi/512
   cos[253]  =  8'b00000001;     //253pi/512
   sin[254]  =  8'b11000000;     //254pi/512
   cos[254]  =  8'b00000000;     //254pi/512
   sin[255]  =  8'b11000000;     //255pi/512
   cos[255]  =  8'b00000000;     //255pi/512
   sin[256]  =  8'b11000000;     //256pi/512
   cos[256]  =  8'b00000000;     //256pi/512
   sin[257]  =  8'b11000000;     //257pi/512
   cos[257]  =  8'b00000000;     //257pi/512
   sin[258]  =  8'b11000000;     //258pi/512
   cos[258]  =  8'b11111111;     //258pi/512
   sin[259]  =  8'b11000000;     //259pi/512
   cos[259]  =  8'b11111111;     //259pi/512
   sin[260]  =  8'b11000000;     //260pi/512
   cos[260]  =  8'b11111110;     //260pi/512
   sin[261]  =  8'b11000000;     //261pi/512
   cos[261]  =  8'b11111110;     //261pi/512
   sin[262]  =  8'b11000000;     //262pi/512
   cos[262]  =  8'b11111110;     //262pi/512
   sin[263]  =  8'b11000000;     //263pi/512
   cos[263]  =  8'b11111101;     //263pi/512
   sin[264]  =  8'b11000000;     //264pi/512
   cos[264]  =  8'b11111101;     //264pi/512
   sin[265]  =  8'b11000000;     //265pi/512
   cos[265]  =  8'b11111100;     //265pi/512
   sin[266]  =  8'b11000000;     //266pi/512
   cos[266]  =  8'b11111100;     //266pi/512
   sin[267]  =  8'b11000000;     //267pi/512
   cos[267]  =  8'b11111100;     //267pi/512
   sin[268]  =  8'b11000000;     //268pi/512
   cos[268]  =  8'b11111011;     //268pi/512
   sin[269]  =  8'b11000000;     //269pi/512
   cos[269]  =  8'b11111011;     //269pi/512
   sin[270]  =  8'b11000000;     //270pi/512
   cos[270]  =  8'b11111011;     //270pi/512
   sin[271]  =  8'b11000000;     //271pi/512
   cos[271]  =  8'b11111010;     //271pi/512
   sin[272]  =  8'b11000000;     //272pi/512
   cos[272]  =  8'b11111010;     //272pi/512
   sin[273]  =  8'b11000000;     //273pi/512
   cos[273]  =  8'b11111001;     //273pi/512
   sin[274]  =  8'b11000000;     //274pi/512
   cos[274]  =  8'b11111001;     //274pi/512
   sin[275]  =  8'b11000000;     //275pi/512
   cos[275]  =  8'b11111001;     //275pi/512
   sin[276]  =  8'b11000000;     //276pi/512
   cos[276]  =  8'b11111000;     //276pi/512
   sin[277]  =  8'b11000001;     //277pi/512
   cos[277]  =  8'b11111000;     //277pi/512
   sin[278]  =  8'b11000001;     //278pi/512
   cos[278]  =  8'b11110111;     //278pi/512
   sin[279]  =  8'b11000001;     //279pi/512
   cos[279]  =  8'b11110111;     //279pi/512
   sin[280]  =  8'b11000001;     //280pi/512
   cos[280]  =  8'b11110111;     //280pi/512
   sin[281]  =  8'b11000001;     //281pi/512
   cos[281]  =  8'b11110110;     //281pi/512
   sin[282]  =  8'b11000001;     //282pi/512
   cos[282]  =  8'b11110110;     //282pi/512
   sin[283]  =  8'b11000001;     //283pi/512
   cos[283]  =  8'b11110101;     //283pi/512
   sin[284]  =  8'b11000001;     //284pi/512
   cos[284]  =  8'b11110101;     //284pi/512
   sin[285]  =  8'b11000001;     //285pi/512
   cos[285]  =  8'b11110101;     //285pi/512
   sin[286]  =  8'b11000001;     //286pi/512
   cos[286]  =  8'b11110100;     //286pi/512
   sin[287]  =  8'b11000001;     //287pi/512
   cos[287]  =  8'b11110100;     //287pi/512
   sin[288]  =  8'b11000001;     //288pi/512
   cos[288]  =  8'b11110100;     //288pi/512
   sin[289]  =  8'b11000001;     //289pi/512
   cos[289]  =  8'b11110011;     //289pi/512
   sin[290]  =  8'b11000001;     //290pi/512
   cos[290]  =  8'b11110011;     //290pi/512
   sin[291]  =  8'b11000001;     //291pi/512
   cos[291]  =  8'b11110010;     //291pi/512
   sin[292]  =  8'b11000010;     //292pi/512
   cos[292]  =  8'b11110010;     //292pi/512
   sin[293]  =  8'b11000010;     //293pi/512
   cos[293]  =  8'b11110010;     //293pi/512
   sin[294]  =  8'b11000010;     //294pi/512
   cos[294]  =  8'b11110001;     //294pi/512
   sin[295]  =  8'b11000010;     //295pi/512
   cos[295]  =  8'b11110001;     //295pi/512
   sin[296]  =  8'b11000010;     //296pi/512
   cos[296]  =  8'b11110000;     //296pi/512
   sin[297]  =  8'b11000010;     //297pi/512
   cos[297]  =  8'b11110000;     //297pi/512
   sin[298]  =  8'b11000010;     //298pi/512
   cos[298]  =  8'b11110000;     //298pi/512
   sin[299]  =  8'b11000010;     //299pi/512
   cos[299]  =  8'b11101111;     //299pi/512
   sin[300]  =  8'b11000010;     //300pi/512
   cos[300]  =  8'b11101111;     //300pi/512
   sin[301]  =  8'b11000010;     //301pi/512
   cos[301]  =  8'b11101111;     //301pi/512
   sin[302]  =  8'b11000011;     //302pi/512
   cos[302]  =  8'b11101110;     //302pi/512
   sin[303]  =  8'b11000011;     //303pi/512
   cos[303]  =  8'b11101110;     //303pi/512
   sin[304]  =  8'b11000011;     //304pi/512
   cos[304]  =  8'b11101101;     //304pi/512
   sin[305]  =  8'b11000011;     //305pi/512
   cos[305]  =  8'b11101101;     //305pi/512
   sin[306]  =  8'b11000011;     //306pi/512
   cos[306]  =  8'b11101101;     //306pi/512
   sin[307]  =  8'b11000011;     //307pi/512
   cos[307]  =  8'b11101100;     //307pi/512
   sin[308]  =  8'b11000011;     //308pi/512
   cos[308]  =  8'b11101100;     //308pi/512
   sin[309]  =  8'b11000011;     //309pi/512
   cos[309]  =  8'b11101100;     //309pi/512
   sin[310]  =  8'b11000011;     //310pi/512
   cos[310]  =  8'b11101011;     //310pi/512
   sin[311]  =  8'b11000100;     //311pi/512
   cos[311]  =  8'b11101011;     //311pi/512
   sin[312]  =  8'b11000100;     //312pi/512
   cos[312]  =  8'b11101010;     //312pi/512
   sin[313]  =  8'b11000100;     //313pi/512
   cos[313]  =  8'b11101010;     //313pi/512
   sin[314]  =  8'b11000100;     //314pi/512
   cos[314]  =  8'b11101010;     //314pi/512
   sin[315]  =  8'b11000100;     //315pi/512
   cos[315]  =  8'b11101001;     //315pi/512
   sin[316]  =  8'b11000100;     //316pi/512
   cos[316]  =  8'b11101001;     //316pi/512
   sin[317]  =  8'b11000100;     //317pi/512
   cos[317]  =  8'b11101001;     //317pi/512
   sin[318]  =  8'b11000101;     //318pi/512
   cos[318]  =  8'b11101000;     //318pi/512
   sin[319]  =  8'b11000101;     //319pi/512
   cos[319]  =  8'b11101000;     //319pi/512
   sin[320]  =  8'b11000101;     //320pi/512
   cos[320]  =  8'b11101000;     //320pi/512
   sin[321]  =  8'b11000101;     //321pi/512
   cos[321]  =  8'b11100111;     //321pi/512
   sin[322]  =  8'b11000101;     //322pi/512
   cos[322]  =  8'b11100111;     //322pi/512
   sin[323]  =  8'b11000101;     //323pi/512
   cos[323]  =  8'b11100110;     //323pi/512
   sin[324]  =  8'b11000101;     //324pi/512
   cos[324]  =  8'b11100110;     //324pi/512
   sin[325]  =  8'b11000110;     //325pi/512
   cos[325]  =  8'b11100110;     //325pi/512
   sin[326]  =  8'b11000110;     //326pi/512
   cos[326]  =  8'b11100101;     //326pi/512
   sin[327]  =  8'b11000110;     //327pi/512
   cos[327]  =  8'b11100101;     //327pi/512
   sin[328]  =  8'b11000110;     //328pi/512
   cos[328]  =  8'b11100101;     //328pi/512
   sin[329]  =  8'b11000110;     //329pi/512
   cos[329]  =  8'b11100100;     //329pi/512
   sin[330]  =  8'b11000110;     //330pi/512
   cos[330]  =  8'b11100100;     //330pi/512
   sin[331]  =  8'b11000111;     //331pi/512
   cos[331]  =  8'b11100100;     //331pi/512
   sin[332]  =  8'b11000111;     //332pi/512
   cos[332]  =  8'b11100011;     //332pi/512
   sin[333]  =  8'b11000111;     //333pi/512
   cos[333]  =  8'b11100011;     //333pi/512
   sin[334]  =  8'b11000111;     //334pi/512
   cos[334]  =  8'b11100011;     //334pi/512
   sin[335]  =  8'b11000111;     //335pi/512
   cos[335]  =  8'b11100010;     //335pi/512
   sin[336]  =  8'b11001000;     //336pi/512
   cos[336]  =  8'b11100010;     //336pi/512
   sin[337]  =  8'b11001000;     //337pi/512
   cos[337]  =  8'b11100001;     //337pi/512
   sin[338]  =  8'b11001000;     //338pi/512
   cos[338]  =  8'b11100001;     //338pi/512
   sin[339]  =  8'b11001000;     //339pi/512
   cos[339]  =  8'b11100001;     //339pi/512
   sin[340]  =  8'b11001000;     //340pi/512
   cos[340]  =  8'b11100000;     //340pi/512
   sin[341]  =  8'b11001001;     //341pi/512
   cos[341]  =  8'b11100000;     //341pi/512
   sin[342]  =  8'b11001001;     //342pi/512
   cos[342]  =  8'b11100000;     //342pi/512
   sin[343]  =  8'b11001001;     //343pi/512
   cos[343]  =  8'b11011111;     //343pi/512
   sin[344]  =  8'b11001001;     //344pi/512
   cos[344]  =  8'b11011111;     //344pi/512
   sin[345]  =  8'b11001001;     //345pi/512
   cos[345]  =  8'b11011111;     //345pi/512
   sin[346]  =  8'b11001010;     //346pi/512
   cos[346]  =  8'b11011110;     //346pi/512
   sin[347]  =  8'b11001010;     //347pi/512
   cos[347]  =  8'b11011110;     //347pi/512
   sin[348]  =  8'b11001010;     //348pi/512
   cos[348]  =  8'b11011110;     //348pi/512
   sin[349]  =  8'b11001010;     //349pi/512
   cos[349]  =  8'b11011101;     //349pi/512
   sin[350]  =  8'b11001010;     //350pi/512
   cos[350]  =  8'b11011101;     //350pi/512
   sin[351]  =  8'b11001011;     //351pi/512
   cos[351]  =  8'b11011101;     //351pi/512
   sin[352]  =  8'b11001011;     //352pi/512
   cos[352]  =  8'b11011100;     //352pi/512
   sin[353]  =  8'b11001011;     //353pi/512
   cos[353]  =  8'b11011100;     //353pi/512
   sin[354]  =  8'b11001011;     //354pi/512
   cos[354]  =  8'b11011100;     //354pi/512
   sin[355]  =  8'b11001011;     //355pi/512
   cos[355]  =  8'b11011011;     //355pi/512
   sin[356]  =  8'b11001100;     //356pi/512
   cos[356]  =  8'b11011011;     //356pi/512
   sin[357]  =  8'b11001100;     //357pi/512
   cos[357]  =  8'b11011011;     //357pi/512
   sin[358]  =  8'b11001100;     //358pi/512
   cos[358]  =  8'b11011011;     //358pi/512
   sin[359]  =  8'b11001100;     //359pi/512
   cos[359]  =  8'b11011010;     //359pi/512
   sin[360]  =  8'b11001101;     //360pi/512
   cos[360]  =  8'b11011010;     //360pi/512
   sin[361]  =  8'b11001101;     //361pi/512
   cos[361]  =  8'b11011010;     //361pi/512
   sin[362]  =  8'b11001101;     //362pi/512
   cos[362]  =  8'b11011001;     //362pi/512
   sin[363]  =  8'b11001101;     //363pi/512
   cos[363]  =  8'b11011001;     //363pi/512
   sin[364]  =  8'b11001110;     //364pi/512
   cos[364]  =  8'b11011001;     //364pi/512
   sin[365]  =  8'b11001110;     //365pi/512
   cos[365]  =  8'b11011000;     //365pi/512
   sin[366]  =  8'b11001110;     //366pi/512
   cos[366]  =  8'b11011000;     //366pi/512
   sin[367]  =  8'b11001110;     //367pi/512
   cos[367]  =  8'b11011000;     //367pi/512
   sin[368]  =  8'b11001111;     //368pi/512
   cos[368]  =  8'b11010111;     //368pi/512
   sin[369]  =  8'b11001111;     //369pi/512
   cos[369]  =  8'b11010111;     //369pi/512
   sin[370]  =  8'b11001111;     //370pi/512
   cos[370]  =  8'b11010111;     //370pi/512
   sin[371]  =  8'b11001111;     //371pi/512
   cos[371]  =  8'b11010110;     //371pi/512
   sin[372]  =  8'b11010000;     //372pi/512
   cos[372]  =  8'b11010110;     //372pi/512
   sin[373]  =  8'b11010000;     //373pi/512
   cos[373]  =  8'b11010110;     //373pi/512
   sin[374]  =  8'b11010000;     //374pi/512
   cos[374]  =  8'b11010110;     //374pi/512
   sin[375]  =  8'b11010000;     //375pi/512
   cos[375]  =  8'b11010101;     //375pi/512
   sin[376]  =  8'b11010001;     //376pi/512
   cos[376]  =  8'b11010101;     //376pi/512
   sin[377]  =  8'b11010001;     //377pi/512
   cos[377]  =  8'b11010101;     //377pi/512
   sin[378]  =  8'b11010001;     //378pi/512
   cos[378]  =  8'b11010100;     //378pi/512
   sin[379]  =  8'b11010001;     //379pi/512
   cos[379]  =  8'b11010100;     //379pi/512
   sin[380]  =  8'b11010010;     //380pi/512
   cos[380]  =  8'b11010100;     //380pi/512
   sin[381]  =  8'b11010010;     //381pi/512
   cos[381]  =  8'b11010100;     //381pi/512
   sin[382]  =  8'b11010010;     //382pi/512
   cos[382]  =  8'b11010011;     //382pi/512
   sin[383]  =  8'b11010010;     //383pi/512
   cos[383]  =  8'b11010011;     //383pi/512
   sin[384]  =  8'b11010011;     //384pi/512
   cos[384]  =  8'b11010011;     //384pi/512
   sin[385]  =  8'b11010011;     //385pi/512
   cos[385]  =  8'b11010010;     //385pi/512
   sin[386]  =  8'b11010011;     //386pi/512
   cos[386]  =  8'b11010010;     //386pi/512
   sin[387]  =  8'b11010100;     //387pi/512
   cos[387]  =  8'b11010010;     //387pi/512
   sin[388]  =  8'b11010100;     //388pi/512
   cos[388]  =  8'b11010010;     //388pi/512
   sin[389]  =  8'b11010100;     //389pi/512
   cos[389]  =  8'b11010001;     //389pi/512
   sin[390]  =  8'b11010100;     //390pi/512
   cos[390]  =  8'b11010001;     //390pi/512
   sin[391]  =  8'b11010101;     //391pi/512
   cos[391]  =  8'b11010001;     //391pi/512
   sin[392]  =  8'b11010101;     //392pi/512
   cos[392]  =  8'b11010001;     //392pi/512
   sin[393]  =  8'b11010101;     //393pi/512
   cos[393]  =  8'b11010000;     //393pi/512
   sin[394]  =  8'b11010110;     //394pi/512
   cos[394]  =  8'b11010000;     //394pi/512
   sin[395]  =  8'b11010110;     //395pi/512
   cos[395]  =  8'b11010000;     //395pi/512
   sin[396]  =  8'b11010110;     //396pi/512
   cos[396]  =  8'b11010000;     //396pi/512
   sin[397]  =  8'b11010110;     //397pi/512
   cos[397]  =  8'b11001111;     //397pi/512
   sin[398]  =  8'b11010111;     //398pi/512
   cos[398]  =  8'b11001111;     //398pi/512
   sin[399]  =  8'b11010111;     //399pi/512
   cos[399]  =  8'b11001111;     //399pi/512
   sin[400]  =  8'b11010111;     //400pi/512
   cos[400]  =  8'b11001111;     //400pi/512
   sin[401]  =  8'b11011000;     //401pi/512
   cos[401]  =  8'b11001110;     //401pi/512
   sin[402]  =  8'b11011000;     //402pi/512
   cos[402]  =  8'b11001110;     //402pi/512
   sin[403]  =  8'b11011000;     //403pi/512
   cos[403]  =  8'b11001110;     //403pi/512
   sin[404]  =  8'b11011001;     //404pi/512
   cos[404]  =  8'b11001110;     //404pi/512
   sin[405]  =  8'b11011001;     //405pi/512
   cos[405]  =  8'b11001101;     //405pi/512
   sin[406]  =  8'b11011001;     //406pi/512
   cos[406]  =  8'b11001101;     //406pi/512
   sin[407]  =  8'b11011010;     //407pi/512
   cos[407]  =  8'b11001101;     //407pi/512
   sin[408]  =  8'b11011010;     //408pi/512
   cos[408]  =  8'b11001101;     //408pi/512
   sin[409]  =  8'b11011010;     //409pi/512
   cos[409]  =  8'b11001100;     //409pi/512
   sin[410]  =  8'b11011011;     //410pi/512
   cos[410]  =  8'b11001100;     //410pi/512
   sin[411]  =  8'b11011011;     //411pi/512
   cos[411]  =  8'b11001100;     //411pi/512
   sin[412]  =  8'b11011011;     //412pi/512
   cos[412]  =  8'b11001100;     //412pi/512
   sin[413]  =  8'b11011011;     //413pi/512
   cos[413]  =  8'b11001011;     //413pi/512
   sin[414]  =  8'b11011100;     //414pi/512
   cos[414]  =  8'b11001011;     //414pi/512
   sin[415]  =  8'b11011100;     //415pi/512
   cos[415]  =  8'b11001011;     //415pi/512
   sin[416]  =  8'b11011100;     //416pi/512
   cos[416]  =  8'b11001011;     //416pi/512
   sin[417]  =  8'b11011101;     //417pi/512
   cos[417]  =  8'b11001011;     //417pi/512
   sin[418]  =  8'b11011101;     //418pi/512
   cos[418]  =  8'b11001010;     //418pi/512
   sin[419]  =  8'b11011101;     //419pi/512
   cos[419]  =  8'b11001010;     //419pi/512
   sin[420]  =  8'b11011110;     //420pi/512
   cos[420]  =  8'b11001010;     //420pi/512
   sin[421]  =  8'b11011110;     //421pi/512
   cos[421]  =  8'b11001010;     //421pi/512
   sin[422]  =  8'b11011110;     //422pi/512
   cos[422]  =  8'b11001010;     //422pi/512
   sin[423]  =  8'b11011111;     //423pi/512
   cos[423]  =  8'b11001001;     //423pi/512
   sin[424]  =  8'b11011111;     //424pi/512
   cos[424]  =  8'b11001001;     //424pi/512
   sin[425]  =  8'b11011111;     //425pi/512
   cos[425]  =  8'b11001001;     //425pi/512
   sin[426]  =  8'b11100000;     //426pi/512
   cos[426]  =  8'b11001001;     //426pi/512
   sin[427]  =  8'b11100000;     //427pi/512
   cos[427]  =  8'b11001001;     //427pi/512
   sin[428]  =  8'b11100000;     //428pi/512
   cos[428]  =  8'b11001000;     //428pi/512
   sin[429]  =  8'b11100001;     //429pi/512
   cos[429]  =  8'b11001000;     //429pi/512
   sin[430]  =  8'b11100001;     //430pi/512
   cos[430]  =  8'b11001000;     //430pi/512
   sin[431]  =  8'b11100001;     //431pi/512
   cos[431]  =  8'b11001000;     //431pi/512
   sin[432]  =  8'b11100010;     //432pi/512
   cos[432]  =  8'b11001000;     //432pi/512
   sin[433]  =  8'b11100010;     //433pi/512
   cos[433]  =  8'b11000111;     //433pi/512
   sin[434]  =  8'b11100011;     //434pi/512
   cos[434]  =  8'b11000111;     //434pi/512
   sin[435]  =  8'b11100011;     //435pi/512
   cos[435]  =  8'b11000111;     //435pi/512
   sin[436]  =  8'b11100011;     //436pi/512
   cos[436]  =  8'b11000111;     //436pi/512
   sin[437]  =  8'b11100100;     //437pi/512
   cos[437]  =  8'b11000111;     //437pi/512
   sin[438]  =  8'b11100100;     //438pi/512
   cos[438]  =  8'b11000110;     //438pi/512
   sin[439]  =  8'b11100100;     //439pi/512
   cos[439]  =  8'b11000110;     //439pi/512
   sin[440]  =  8'b11100101;     //440pi/512
   cos[440]  =  8'b11000110;     //440pi/512
   sin[441]  =  8'b11100101;     //441pi/512
   cos[441]  =  8'b11000110;     //441pi/512
   sin[442]  =  8'b11100101;     //442pi/512
   cos[442]  =  8'b11000110;     //442pi/512
   sin[443]  =  8'b11100110;     //443pi/512
   cos[443]  =  8'b11000110;     //443pi/512
   sin[444]  =  8'b11100110;     //444pi/512
   cos[444]  =  8'b11000101;     //444pi/512
   sin[445]  =  8'b11100110;     //445pi/512
   cos[445]  =  8'b11000101;     //445pi/512
   sin[446]  =  8'b11100111;     //446pi/512
   cos[446]  =  8'b11000101;     //446pi/512
   sin[447]  =  8'b11100111;     //447pi/512
   cos[447]  =  8'b11000101;     //447pi/512
   sin[448]  =  8'b11101000;     //448pi/512
   cos[448]  =  8'b11000101;     //448pi/512
   sin[449]  =  8'b11101000;     //449pi/512
   cos[449]  =  8'b11000101;     //449pi/512
   sin[450]  =  8'b11101000;     //450pi/512
   cos[450]  =  8'b11000101;     //450pi/512
   sin[451]  =  8'b11101001;     //451pi/512
   cos[451]  =  8'b11000100;     //451pi/512
   sin[452]  =  8'b11101001;     //452pi/512
   cos[452]  =  8'b11000100;     //452pi/512
   sin[453]  =  8'b11101001;     //453pi/512
   cos[453]  =  8'b11000100;     //453pi/512
   sin[454]  =  8'b11101010;     //454pi/512
   cos[454]  =  8'b11000100;     //454pi/512
   sin[455]  =  8'b11101010;     //455pi/512
   cos[455]  =  8'b11000100;     //455pi/512
   sin[456]  =  8'b11101010;     //456pi/512
   cos[456]  =  8'b11000100;     //456pi/512
   sin[457]  =  8'b11101011;     //457pi/512
   cos[457]  =  8'b11000100;     //457pi/512
   sin[458]  =  8'b11101011;     //458pi/512
   cos[458]  =  8'b11000011;     //458pi/512
   sin[459]  =  8'b11101100;     //459pi/512
   cos[459]  =  8'b11000011;     //459pi/512
   sin[460]  =  8'b11101100;     //460pi/512
   cos[460]  =  8'b11000011;     //460pi/512
   sin[461]  =  8'b11101100;     //461pi/512
   cos[461]  =  8'b11000011;     //461pi/512
   sin[462]  =  8'b11101101;     //462pi/512
   cos[462]  =  8'b11000011;     //462pi/512
   sin[463]  =  8'b11101101;     //463pi/512
   cos[463]  =  8'b11000011;     //463pi/512
   sin[464]  =  8'b11101101;     //464pi/512
   cos[464]  =  8'b11000011;     //464pi/512
   sin[465]  =  8'b11101110;     //465pi/512
   cos[465]  =  8'b11000011;     //465pi/512
   sin[466]  =  8'b11101110;     //466pi/512
   cos[466]  =  8'b11000011;     //466pi/512
   sin[467]  =  8'b11101111;     //467pi/512
   cos[467]  =  8'b11000010;     //467pi/512
   sin[468]  =  8'b11101111;     //468pi/512
   cos[468]  =  8'b11000010;     //468pi/512
   sin[469]  =  8'b11101111;     //469pi/512
   cos[469]  =  8'b11000010;     //469pi/512
   sin[470]  =  8'b11110000;     //470pi/512
   cos[470]  =  8'b11000010;     //470pi/512
   sin[471]  =  8'b11110000;     //471pi/512
   cos[471]  =  8'b11000010;     //471pi/512
   sin[472]  =  8'b11110000;     //472pi/512
   cos[472]  =  8'b11000010;     //472pi/512
   sin[473]  =  8'b11110001;     //473pi/512
   cos[473]  =  8'b11000010;     //473pi/512
   sin[474]  =  8'b11110001;     //474pi/512
   cos[474]  =  8'b11000010;     //474pi/512
   sin[475]  =  8'b11110010;     //475pi/512
   cos[475]  =  8'b11000010;     //475pi/512
   sin[476]  =  8'b11110010;     //476pi/512
   cos[476]  =  8'b11000010;     //476pi/512
   sin[477]  =  8'b11110010;     //477pi/512
   cos[477]  =  8'b11000001;     //477pi/512
   sin[478]  =  8'b11110011;     //478pi/512
   cos[478]  =  8'b11000001;     //478pi/512
   sin[479]  =  8'b11110011;     //479pi/512
   cos[479]  =  8'b11000001;     //479pi/512
   sin[480]  =  8'b11110100;     //480pi/512
   cos[480]  =  8'b11000001;     //480pi/512
   sin[481]  =  8'b11110100;     //481pi/512
   cos[481]  =  8'b11000001;     //481pi/512
   sin[482]  =  8'b11110100;     //482pi/512
   cos[482]  =  8'b11000001;     //482pi/512
   sin[483]  =  8'b11110101;     //483pi/512
   cos[483]  =  8'b11000001;     //483pi/512
   sin[484]  =  8'b11110101;     //484pi/512
   cos[484]  =  8'b11000001;     //484pi/512
   sin[485]  =  8'b11110101;     //485pi/512
   cos[485]  =  8'b11000001;     //485pi/512
   sin[486]  =  8'b11110110;     //486pi/512
   cos[486]  =  8'b11000001;     //486pi/512
   sin[487]  =  8'b11110110;     //487pi/512
   cos[487]  =  8'b11000001;     //487pi/512
   sin[488]  =  8'b11110111;     //488pi/512
   cos[488]  =  8'b11000001;     //488pi/512
   sin[489]  =  8'b11110111;     //489pi/512
   cos[489]  =  8'b11000001;     //489pi/512
   sin[490]  =  8'b11110111;     //490pi/512
   cos[490]  =  8'b11000001;     //490pi/512
   sin[491]  =  8'b11111000;     //491pi/512
   cos[491]  =  8'b11000001;     //491pi/512
   sin[492]  =  8'b11111000;     //492pi/512
   cos[492]  =  8'b11000000;     //492pi/512
   sin[493]  =  8'b11111001;     //493pi/512
   cos[493]  =  8'b11000000;     //493pi/512
   sin[494]  =  8'b11111001;     //494pi/512
   cos[494]  =  8'b11000000;     //494pi/512
   sin[495]  =  8'b11111001;     //495pi/512
   cos[495]  =  8'b11000000;     //495pi/512
   sin[496]  =  8'b11111010;     //496pi/512
   cos[496]  =  8'b11000000;     //496pi/512
   sin[497]  =  8'b11111010;     //497pi/512
   cos[497]  =  8'b11000000;     //497pi/512
   sin[498]  =  8'b11111011;     //498pi/512
   cos[498]  =  8'b11000000;     //498pi/512
   sin[499]  =  8'b11111011;     //499pi/512
   cos[499]  =  8'b11000000;     //499pi/512
   sin[500]  =  8'b11111011;     //500pi/512
   cos[500]  =  8'b11000000;     //500pi/512
   sin[501]  =  8'b11111100;     //501pi/512
   cos[501]  =  8'b11000000;     //501pi/512
   sin[502]  =  8'b11111100;     //502pi/512
   cos[502]  =  8'b11000000;     //502pi/512
   sin[503]  =  8'b11111100;     //503pi/512
   cos[503]  =  8'b11000000;     //503pi/512
   sin[504]  =  8'b11111101;     //504pi/512
   cos[504]  =  8'b11000000;     //504pi/512
   sin[505]  =  8'b11111101;     //505pi/512
   cos[505]  =  8'b11000000;     //505pi/512
   sin[506]  =  8'b11111110;     //506pi/512
   cos[506]  =  8'b11000000;     //506pi/512
   sin[507]  =  8'b11111110;     //507pi/512
   cos[507]  =  8'b11000000;     //507pi/512
   sin[508]  =  8'b11111110;     //508pi/512
   cos[508]  =  8'b11000000;     //508pi/512
   sin[509]  =  8'b11111111;     //509pi/512
   cos[509]  =  8'b11000000;     //509pi/512
   sin[510]  =  8'b11111111;     //510pi/512
   cos[510]  =  8'b11000000;     //510pi/512
   sin[511]  =  8'b00000000;     //511pi/512
   cos[511]  =  8'b11000000;     //511pi/512
/////////////////////////////////////////////////////////////////

   m_sin[0]  =  8'b00000000;     //0pi/512
   m_cos[0]  =  8'b01000000;     //0pi/512
   m_sin[1]  =  8'b00000000;     //1pi/512
   m_cos[1]  =  8'b00111111;     //1pi/512
   m_sin[2]  =  8'b11111111;     //2pi/512
   m_cos[2]  =  8'b00111111;     //2pi/512
   m_sin[3]  =  8'b11111111;     //3pi/512
   m_cos[3]  =  8'b00111111;     //3pi/512
   m_sin[4]  =  8'b11111111;     //4pi/512
   m_cos[4]  =  8'b00111111;     //4pi/512
   m_sin[5]  =  8'b11111110;     //5pi/512
   m_cos[5]  =  8'b00111111;     //5pi/512
   m_sin[6]  =  8'b11111110;     //6pi/512
   m_cos[6]  =  8'b00111111;     //6pi/512
   m_sin[7]  =  8'b11111110;     //7pi/512
   m_cos[7]  =  8'b00111111;     //7pi/512
   m_sin[8]  =  8'b11111101;     //8pi/512
   m_cos[8]  =  8'b00111111;     //8pi/512
   m_sin[9]  =  8'b11111101;     //9pi/512
   m_cos[9]  =  8'b00111111;     //9pi/512
   m_sin[10]  =  8'b11111101;     //10pi/512
   m_cos[10]  =  8'b00111111;     //10pi/512
   m_sin[11]  =  8'b11111101;     //11pi/512
   m_cos[11]  =  8'b00111111;     //11pi/512
   m_sin[12]  =  8'b11111100;     //12pi/512
   m_cos[12]  =  8'b00111111;     //12pi/512
   m_sin[13]  =  8'b11111100;     //13pi/512
   m_cos[13]  =  8'b00111111;     //13pi/512
   m_sin[14]  =  8'b11111100;     //14pi/512
   m_cos[14]  =  8'b00111111;     //14pi/512
   m_sin[15]  =  8'b11111011;     //15pi/512
   m_cos[15]  =  8'b00111111;     //15pi/512
   m_sin[16]  =  8'b11111011;     //16pi/512
   m_cos[16]  =  8'b00111111;     //16pi/512
   m_sin[17]  =  8'b11111011;     //17pi/512
   m_cos[17]  =  8'b00111111;     //17pi/512
   m_sin[18]  =  8'b11111010;     //18pi/512
   m_cos[18]  =  8'b00111111;     //18pi/512
   m_sin[19]  =  8'b11111010;     //19pi/512
   m_cos[19]  =  8'b00111111;     //19pi/512
   m_sin[20]  =  8'b11111010;     //20pi/512
   m_cos[20]  =  8'b00111111;     //20pi/512
   m_sin[21]  =  8'b11111001;     //21pi/512
   m_cos[21]  =  8'b00111111;     //21pi/512
   m_sin[22]  =  8'b11111001;     //22pi/512
   m_cos[22]  =  8'b00111111;     //22pi/512
   m_sin[23]  =  8'b11111001;     //23pi/512
   m_cos[23]  =  8'b00111111;     //23pi/512
   m_sin[24]  =  8'b11111000;     //24pi/512
   m_cos[24]  =  8'b00111111;     //24pi/512
   m_sin[25]  =  8'b11111000;     //25pi/512
   m_cos[25]  =  8'b00111111;     //25pi/512
   m_sin[26]  =  8'b11111000;     //26pi/512
   m_cos[26]  =  8'b00111111;     //26pi/512
   m_sin[27]  =  8'b11111000;     //27pi/512
   m_cos[27]  =  8'b00111111;     //27pi/512
   m_sin[28]  =  8'b11110111;     //28pi/512
   m_cos[28]  =  8'b00111111;     //28pi/512
   m_sin[29]  =  8'b11110111;     //29pi/512
   m_cos[29]  =  8'b00111111;     //29pi/512
   m_sin[30]  =  8'b11110111;     //30pi/512
   m_cos[30]  =  8'b00111111;     //30pi/512
   m_sin[31]  =  8'b11110110;     //31pi/512
   m_cos[31]  =  8'b00111111;     //31pi/512
   m_sin[32]  =  8'b11110110;     //32pi/512
   m_cos[32]  =  8'b00111111;     //32pi/512
   m_sin[33]  =  8'b11110110;     //33pi/512
   m_cos[33]  =  8'b00111111;     //33pi/512
   m_sin[34]  =  8'b11110101;     //34pi/512
   m_cos[34]  =  8'b00111111;     //34pi/512
   m_sin[35]  =  8'b11110101;     //35pi/512
   m_cos[35]  =  8'b00111111;     //35pi/512
   m_sin[36]  =  8'b11110101;     //36pi/512
   m_cos[36]  =  8'b00111111;     //36pi/512
   m_sin[37]  =  8'b11110100;     //37pi/512
   m_cos[37]  =  8'b00111110;     //37pi/512
   m_sin[38]  =  8'b11110100;     //38pi/512
   m_cos[38]  =  8'b00111110;     //38pi/512
   m_sin[39]  =  8'b11110100;     //39pi/512
   m_cos[39]  =  8'b00111110;     //39pi/512
   m_sin[40]  =  8'b11110100;     //40pi/512
   m_cos[40]  =  8'b00111110;     //40pi/512
   m_sin[41]  =  8'b11110011;     //41pi/512
   m_cos[41]  =  8'b00111110;     //41pi/512
   m_sin[42]  =  8'b11110011;     //42pi/512
   m_cos[42]  =  8'b00111110;     //42pi/512
   m_sin[43]  =  8'b11110011;     //43pi/512
   m_cos[43]  =  8'b00111110;     //43pi/512
   m_sin[44]  =  8'b11110010;     //44pi/512
   m_cos[44]  =  8'b00111110;     //44pi/512
   m_sin[45]  =  8'b11110010;     //45pi/512
   m_cos[45]  =  8'b00111110;     //45pi/512
   m_sin[46]  =  8'b11110010;     //46pi/512
   m_cos[46]  =  8'b00111110;     //46pi/512
   m_sin[47]  =  8'b11110001;     //47pi/512
   m_cos[47]  =  8'b00111110;     //47pi/512
   m_sin[48]  =  8'b11110001;     //48pi/512
   m_cos[48]  =  8'b00111110;     //48pi/512
   m_sin[49]  =  8'b11110001;     //49pi/512
   m_cos[49]  =  8'b00111110;     //49pi/512
   m_sin[50]  =  8'b11110000;     //50pi/512
   m_cos[50]  =  8'b00111110;     //50pi/512
   m_sin[51]  =  8'b11110000;     //51pi/512
   m_cos[51]  =  8'b00111110;     //51pi/512
   m_sin[52]  =  8'b11110000;     //52pi/512
   m_cos[52]  =  8'b00111101;     //52pi/512
   m_sin[53]  =  8'b11110000;     //53pi/512
   m_cos[53]  =  8'b00111101;     //53pi/512
   m_sin[54]  =  8'b11101111;     //54pi/512
   m_cos[54]  =  8'b00111101;     //54pi/512
   m_sin[55]  =  8'b11101111;     //55pi/512
   m_cos[55]  =  8'b00111101;     //55pi/512
   m_sin[56]  =  8'b11101111;     //56pi/512
   m_cos[56]  =  8'b00111101;     //56pi/512
   m_sin[57]  =  8'b11101110;     //57pi/512
   m_cos[57]  =  8'b00111101;     //57pi/512
   m_sin[58]  =  8'b11101110;     //58pi/512
   m_cos[58]  =  8'b00111101;     //58pi/512
   m_sin[59]  =  8'b11101110;     //59pi/512
   m_cos[59]  =  8'b00111101;     //59pi/512
   m_sin[60]  =  8'b11101101;     //60pi/512
   m_cos[60]  =  8'b00111101;     //60pi/512
   m_sin[61]  =  8'b11101101;     //61pi/512
   m_cos[61]  =  8'b00111101;     //61pi/512
   m_sin[62]  =  8'b11101101;     //62pi/512
   m_cos[62]  =  8'b00111101;     //62pi/512
   m_sin[63]  =  8'b11101101;     //63pi/512
   m_cos[63]  =  8'b00111100;     //63pi/512
   m_sin[64]  =  8'b11101100;     //64pi/512
   m_cos[64]  =  8'b00111100;     //64pi/512
   m_sin[65]  =  8'b11101100;     //65pi/512
   m_cos[65]  =  8'b00111100;     //65pi/512
   m_sin[66]  =  8'b11101100;     //66pi/512
   m_cos[66]  =  8'b00111100;     //66pi/512
   m_sin[67]  =  8'b11101011;     //67pi/512
   m_cos[67]  =  8'b00111100;     //67pi/512
   m_sin[68]  =  8'b11101011;     //68pi/512
   m_cos[68]  =  8'b00111100;     //68pi/512
   m_sin[69]  =  8'b11101011;     //69pi/512
   m_cos[69]  =  8'b00111100;     //69pi/512
   m_sin[70]  =  8'b11101010;     //70pi/512
   m_cos[70]  =  8'b00111100;     //70pi/512
   m_sin[71]  =  8'b11101010;     //71pi/512
   m_cos[71]  =  8'b00111100;     //71pi/512
   m_sin[72]  =  8'b11101010;     //72pi/512
   m_cos[72]  =  8'b00111100;     //72pi/512
   m_sin[73]  =  8'b11101010;     //73pi/512
   m_cos[73]  =  8'b00111011;     //73pi/512
   m_sin[74]  =  8'b11101001;     //74pi/512
   m_cos[74]  =  8'b00111011;     //74pi/512
   m_sin[75]  =  8'b11101001;     //75pi/512
   m_cos[75]  =  8'b00111011;     //75pi/512
   m_sin[76]  =  8'b11101001;     //76pi/512
   m_cos[76]  =  8'b00111011;     //76pi/512
   m_sin[77]  =  8'b11101000;     //77pi/512
   m_cos[77]  =  8'b00111011;     //77pi/512
   m_sin[78]  =  8'b11101000;     //78pi/512
   m_cos[78]  =  8'b00111011;     //78pi/512
   m_sin[79]  =  8'b11101000;     //79pi/512
   m_cos[79]  =  8'b00111011;     //79pi/512
   m_sin[80]  =  8'b11101000;     //80pi/512
   m_cos[80]  =  8'b00111011;     //80pi/512
   m_sin[81]  =  8'b11100111;     //81pi/512
   m_cos[81]  =  8'b00111011;     //81pi/512
   m_sin[82]  =  8'b11100111;     //82pi/512
   m_cos[82]  =  8'b00111010;     //82pi/512
   m_sin[83]  =  8'b11100111;     //83pi/512
   m_cos[83]  =  8'b00111010;     //83pi/512
   m_sin[84]  =  8'b11100110;     //84pi/512
   m_cos[84]  =  8'b00111010;     //84pi/512
   m_sin[85]  =  8'b11100110;     //85pi/512
   m_cos[85]  =  8'b00111010;     //85pi/512
   m_sin[86]  =  8'b11100110;     //86pi/512
   m_cos[86]  =  8'b00111010;     //86pi/512
   m_sin[87]  =  8'b11100101;     //87pi/512
   m_cos[87]  =  8'b00111010;     //87pi/512
   m_sin[88]  =  8'b11100101;     //88pi/512
   m_cos[88]  =  8'b00111010;     //88pi/512
   m_sin[89]  =  8'b11100101;     //89pi/512
   m_cos[89]  =  8'b00111001;     //89pi/512
   m_sin[90]  =  8'b11100101;     //90pi/512
   m_cos[90]  =  8'b00111001;     //90pi/512
   m_sin[91]  =  8'b11100100;     //91pi/512
   m_cos[91]  =  8'b00111001;     //91pi/512
   m_sin[92]  =  8'b11100100;     //92pi/512
   m_cos[92]  =  8'b00111001;     //92pi/512
   m_sin[93]  =  8'b11100100;     //93pi/512
   m_cos[93]  =  8'b00111001;     //93pi/512
   m_sin[94]  =  8'b11100100;     //94pi/512
   m_cos[94]  =  8'b00111001;     //94pi/512
   m_sin[95]  =  8'b11100011;     //95pi/512
   m_cos[95]  =  8'b00111001;     //95pi/512
   m_sin[96]  =  8'b11100011;     //96pi/512
   m_cos[96]  =  8'b00111001;     //96pi/512
   m_sin[97]  =  8'b11100011;     //97pi/512
   m_cos[97]  =  8'b00111000;     //97pi/512
   m_sin[98]  =  8'b11100010;     //98pi/512
   m_cos[98]  =  8'b00111000;     //98pi/512
   m_sin[99]  =  8'b11100010;     //99pi/512
   m_cos[99]  =  8'b00111000;     //99pi/512
   m_sin[100]  =  8'b11100010;     //100pi/512
   m_cos[100]  =  8'b00111000;     //100pi/512
   m_sin[101]  =  8'b11100010;     //101pi/512
   m_cos[101]  =  8'b00111000;     //101pi/512
   m_sin[102]  =  8'b11100001;     //102pi/512
   m_cos[102]  =  8'b00111000;     //102pi/512
   m_sin[103]  =  8'b11100001;     //103pi/512
   m_cos[103]  =  8'b00110111;     //103pi/512
   m_sin[104]  =  8'b11100001;     //104pi/512
   m_cos[104]  =  8'b00110111;     //104pi/512
   m_sin[105]  =  8'b11100000;     //105pi/512
   m_cos[105]  =  8'b00110111;     //105pi/512
   m_sin[106]  =  8'b11100000;     //106pi/512
   m_cos[106]  =  8'b00110111;     //106pi/512
   m_sin[107]  =  8'b11100000;     //107pi/512
   m_cos[107]  =  8'b00110111;     //107pi/512
   m_sin[108]  =  8'b11100000;     //108pi/512
   m_cos[108]  =  8'b00110111;     //108pi/512
   m_sin[109]  =  8'b11011111;     //109pi/512
   m_cos[109]  =  8'b00110111;     //109pi/512
   m_sin[110]  =  8'b11011111;     //110pi/512
   m_cos[110]  =  8'b00110110;     //110pi/512
   m_sin[111]  =  8'b11011111;     //111pi/512
   m_cos[111]  =  8'b00110110;     //111pi/512
   m_sin[112]  =  8'b11011111;     //112pi/512
   m_cos[112]  =  8'b00110110;     //112pi/512
   m_sin[113]  =  8'b11011110;     //113pi/512
   m_cos[113]  =  8'b00110110;     //113pi/512
   m_sin[114]  =  8'b11011110;     //114pi/512
   m_cos[114]  =  8'b00110110;     //114pi/512
   m_sin[115]  =  8'b11011110;     //115pi/512
   m_cos[115]  =  8'b00110110;     //115pi/512
   m_sin[116]  =  8'b11011101;     //116pi/512
   m_cos[116]  =  8'b00110101;     //116pi/512
   m_sin[117]  =  8'b11011101;     //117pi/512
   m_cos[117]  =  8'b00110101;     //117pi/512
   m_sin[118]  =  8'b11011101;     //118pi/512
   m_cos[118]  =  8'b00110101;     //118pi/512
   m_sin[119]  =  8'b11011101;     //119pi/512
   m_cos[119]  =  8'b00110101;     //119pi/512
   m_sin[120]  =  8'b11011100;     //120pi/512
   m_cos[120]  =  8'b00110101;     //120pi/512
   m_sin[121]  =  8'b11011100;     //121pi/512
   m_cos[121]  =  8'b00110101;     //121pi/512
   m_sin[122]  =  8'b11011100;     //122pi/512
   m_cos[122]  =  8'b00110100;     //122pi/512
   m_sin[123]  =  8'b11011100;     //123pi/512
   m_cos[123]  =  8'b00110100;     //123pi/512
   m_sin[124]  =  8'b11011011;     //124pi/512
   m_cos[124]  =  8'b00110100;     //124pi/512
   m_sin[125]  =  8'b11011011;     //125pi/512
   m_cos[125]  =  8'b00110100;     //125pi/512
   m_sin[126]  =  8'b11011011;     //126pi/512
   m_cos[126]  =  8'b00110100;     //126pi/512
   m_sin[127]  =  8'b11011011;     //127pi/512
   m_cos[127]  =  8'b00110011;     //127pi/512
   m_sin[128]  =  8'b11011010;     //128pi/512
   m_cos[128]  =  8'b00110011;     //128pi/512
   m_sin[129]  =  8'b11011010;     //129pi/512
   m_cos[129]  =  8'b00110011;     //129pi/512
   m_sin[130]  =  8'b11011010;     //130pi/512
   m_cos[130]  =  8'b00110011;     //130pi/512
   m_sin[131]  =  8'b11011010;     //131pi/512
   m_cos[131]  =  8'b00110011;     //131pi/512
   m_sin[132]  =  8'b11011001;     //132pi/512
   m_cos[132]  =  8'b00110011;     //132pi/512
   m_sin[133]  =  8'b11011001;     //133pi/512
   m_cos[133]  =  8'b00110010;     //133pi/512
   m_sin[134]  =  8'b11011001;     //134pi/512
   m_cos[134]  =  8'b00110010;     //134pi/512
   m_sin[135]  =  8'b11011001;     //135pi/512
   m_cos[135]  =  8'b00110010;     //135pi/512
   m_sin[136]  =  8'b11011000;     //136pi/512
   m_cos[136]  =  8'b00110010;     //136pi/512
   m_sin[137]  =  8'b11011000;     //137pi/512
   m_cos[137]  =  8'b00110010;     //137pi/512
   m_sin[138]  =  8'b11011000;     //138pi/512
   m_cos[138]  =  8'b00110001;     //138pi/512
   m_sin[139]  =  8'b11011000;     //139pi/512
   m_cos[139]  =  8'b00110001;     //139pi/512
   m_sin[140]  =  8'b11010111;     //140pi/512
   m_cos[140]  =  8'b00110001;     //140pi/512
   m_sin[141]  =  8'b11010111;     //141pi/512
   m_cos[141]  =  8'b00110001;     //141pi/512
   m_sin[142]  =  8'b11010111;     //142pi/512
   m_cos[142]  =  8'b00110001;     //142pi/512
   m_sin[143]  =  8'b11010111;     //143pi/512
   m_cos[143]  =  8'b00110000;     //143pi/512
   m_sin[144]  =  8'b11010110;     //144pi/512
   m_cos[144]  =  8'b00110000;     //144pi/512
   m_sin[145]  =  8'b11010110;     //145pi/512
   m_cos[145]  =  8'b00110000;     //145pi/512
   m_sin[146]  =  8'b11010110;     //146pi/512
   m_cos[146]  =  8'b00110000;     //146pi/512
   m_sin[147]  =  8'b11010110;     //147pi/512
   m_cos[147]  =  8'b00110000;     //147pi/512
   m_sin[148]  =  8'b11010101;     //148pi/512
   m_cos[148]  =  8'b00101111;     //148pi/512
   m_sin[149]  =  8'b11010101;     //149pi/512
   m_cos[149]  =  8'b00101111;     //149pi/512
   m_sin[150]  =  8'b11010101;     //150pi/512
   m_cos[150]  =  8'b00101111;     //150pi/512
   m_sin[151]  =  8'b11010101;     //151pi/512
   m_cos[151]  =  8'b00101111;     //151pi/512
   m_sin[152]  =  8'b11010101;     //152pi/512
   m_cos[152]  =  8'b00101110;     //152pi/512
   m_sin[153]  =  8'b11010100;     //153pi/512
   m_cos[153]  =  8'b00101110;     //153pi/512
   m_sin[154]  =  8'b11010100;     //154pi/512
   m_cos[154]  =  8'b00101110;     //154pi/512
   m_sin[155]  =  8'b11010100;     //155pi/512
   m_cos[155]  =  8'b00101110;     //155pi/512
   m_sin[156]  =  8'b11010100;     //156pi/512
   m_cos[156]  =  8'b00101110;     //156pi/512
   m_sin[157]  =  8'b11010011;     //157pi/512
   m_cos[157]  =  8'b00101101;     //157pi/512
   m_sin[158]  =  8'b11010011;     //158pi/512
   m_cos[158]  =  8'b00101101;     //158pi/512
   m_sin[159]  =  8'b11010011;     //159pi/512
   m_cos[159]  =  8'b00101101;     //159pi/512
   m_sin[160]  =  8'b11010011;     //160pi/512
   m_cos[160]  =  8'b00101101;     //160pi/512
   m_sin[161]  =  8'b11010011;     //161pi/512
   m_cos[161]  =  8'b00101101;     //161pi/512
   m_sin[162]  =  8'b11010010;     //162pi/512
   m_cos[162]  =  8'b00101100;     //162pi/512
   m_sin[163]  =  8'b11010010;     //163pi/512
   m_cos[163]  =  8'b00101100;     //163pi/512
   m_sin[164]  =  8'b11010010;     //164pi/512
   m_cos[164]  =  8'b00101100;     //164pi/512
   m_sin[165]  =  8'b11010010;     //165pi/512
   m_cos[165]  =  8'b00101100;     //165pi/512
   m_sin[166]  =  8'b11010001;     //166pi/512
   m_cos[166]  =  8'b00101011;     //166pi/512
   m_sin[167]  =  8'b11010001;     //167pi/512
   m_cos[167]  =  8'b00101011;     //167pi/512
   m_sin[168]  =  8'b11010001;     //168pi/512
   m_cos[168]  =  8'b00101011;     //168pi/512
   m_sin[169]  =  8'b11010001;     //169pi/512
   m_cos[169]  =  8'b00101011;     //169pi/512
   m_sin[170]  =  8'b11010001;     //170pi/512
   m_cos[170]  =  8'b00101010;     //170pi/512
   m_sin[171]  =  8'b11010000;     //171pi/512
   m_cos[171]  =  8'b00101010;     //171pi/512
   m_sin[172]  =  8'b11010000;     //172pi/512
   m_cos[172]  =  8'b00101010;     //172pi/512
   m_sin[173]  =  8'b11010000;     //173pi/512
   m_cos[173]  =  8'b00101010;     //173pi/512
   m_sin[174]  =  8'b11010000;     //174pi/512
   m_cos[174]  =  8'b00101010;     //174pi/512
   m_sin[175]  =  8'b11010000;     //175pi/512
   m_cos[175]  =  8'b00101001;     //175pi/512
   m_sin[176]  =  8'b11001111;     //176pi/512
   m_cos[176]  =  8'b00101001;     //176pi/512
   m_sin[177]  =  8'b11001111;     //177pi/512
   m_cos[177]  =  8'b00101001;     //177pi/512
   m_sin[178]  =  8'b11001111;     //178pi/512
   m_cos[178]  =  8'b00101001;     //178pi/512
   m_sin[179]  =  8'b11001111;     //179pi/512
   m_cos[179]  =  8'b00101000;     //179pi/512
   m_sin[180]  =  8'b11001111;     //180pi/512
   m_cos[180]  =  8'b00101000;     //180pi/512
   m_sin[181]  =  8'b11001110;     //181pi/512
   m_cos[181]  =  8'b00101000;     //181pi/512
   m_sin[182]  =  8'b11001110;     //182pi/512
   m_cos[182]  =  8'b00101000;     //182pi/512
   m_sin[183]  =  8'b11001110;     //183pi/512
   m_cos[183]  =  8'b00100111;     //183pi/512
   m_sin[184]  =  8'b11001110;     //184pi/512
   m_cos[184]  =  8'b00100111;     //184pi/512
   m_sin[185]  =  8'b11001110;     //185pi/512
   m_cos[185]  =  8'b00100111;     //185pi/512
   m_sin[186]  =  8'b11001101;     //186pi/512
   m_cos[186]  =  8'b00100111;     //186pi/512
   m_sin[187]  =  8'b11001101;     //187pi/512
   m_cos[187]  =  8'b00100110;     //187pi/512
   m_sin[188]  =  8'b11001101;     //188pi/512
   m_cos[188]  =  8'b00100110;     //188pi/512
   m_sin[189]  =  8'b11001101;     //189pi/512
   m_cos[189]  =  8'b00100110;     //189pi/512
   m_sin[190]  =  8'b11001101;     //190pi/512
   m_cos[190]  =  8'b00100110;     //190pi/512
   m_sin[191]  =  8'b11001100;     //191pi/512
   m_cos[191]  =  8'b00100101;     //191pi/512
   m_sin[192]  =  8'b11001100;     //192pi/512
   m_cos[192]  =  8'b00100101;     //192pi/512
   m_sin[193]  =  8'b11001100;     //193pi/512
   m_cos[193]  =  8'b00100101;     //193pi/512
   m_sin[194]  =  8'b11001100;     //194pi/512
   m_cos[194]  =  8'b00100101;     //194pi/512
   m_sin[195]  =  8'b11001100;     //195pi/512
   m_cos[195]  =  8'b00100100;     //195pi/512
   m_sin[196]  =  8'b11001011;     //196pi/512
   m_cos[196]  =  8'b00100100;     //196pi/512
   m_sin[197]  =  8'b11001011;     //197pi/512
   m_cos[197]  =  8'b00100100;     //197pi/512
   m_sin[198]  =  8'b11001011;     //198pi/512
   m_cos[198]  =  8'b00100100;     //198pi/512
   m_sin[199]  =  8'b11001011;     //199pi/512
   m_cos[199]  =  8'b00100011;     //199pi/512
   m_sin[200]  =  8'b11001011;     //200pi/512
   m_cos[200]  =  8'b00100011;     //200pi/512
   m_sin[201]  =  8'b11001011;     //201pi/512
   m_cos[201]  =  8'b00100011;     //201pi/512
   m_sin[202]  =  8'b11001010;     //202pi/512
   m_cos[202]  =  8'b00100011;     //202pi/512
   m_sin[203]  =  8'b11001010;     //203pi/512
   m_cos[203]  =  8'b00100010;     //203pi/512
   m_sin[204]  =  8'b11001010;     //204pi/512
   m_cos[204]  =  8'b00100010;     //204pi/512
   m_sin[205]  =  8'b11001010;     //205pi/512
   m_cos[205]  =  8'b00100010;     //205pi/512
   m_sin[206]  =  8'b11001010;     //206pi/512
   m_cos[206]  =  8'b00100001;     //206pi/512
   m_sin[207]  =  8'b11001010;     //207pi/512
   m_cos[207]  =  8'b00100001;     //207pi/512
   m_sin[208]  =  8'b11001001;     //208pi/512
   m_cos[208]  =  8'b00100001;     //208pi/512
   m_sin[209]  =  8'b11001001;     //209pi/512
   m_cos[209]  =  8'b00100001;     //209pi/512
   m_sin[210]  =  8'b11001001;     //210pi/512
   m_cos[210]  =  8'b00100000;     //210pi/512
   m_sin[211]  =  8'b11001001;     //211pi/512
   m_cos[211]  =  8'b00100000;     //211pi/512
   m_sin[212]  =  8'b11001001;     //212pi/512
   m_cos[212]  =  8'b00100000;     //212pi/512
   m_sin[213]  =  8'b11001001;     //213pi/512
   m_cos[213]  =  8'b00100000;     //213pi/512
   m_sin[214]  =  8'b11001000;     //214pi/512
   m_cos[214]  =  8'b00011111;     //214pi/512
   m_sin[215]  =  8'b11001000;     //215pi/512
   m_cos[215]  =  8'b00011111;     //215pi/512
   m_sin[216]  =  8'b11001000;     //216pi/512
   m_cos[216]  =  8'b00011111;     //216pi/512
   m_sin[217]  =  8'b11001000;     //217pi/512
   m_cos[217]  =  8'b00011110;     //217pi/512
   m_sin[218]  =  8'b11001000;     //218pi/512
   m_cos[218]  =  8'b00011110;     //218pi/512
   m_sin[219]  =  8'b11001000;     //219pi/512
   m_cos[219]  =  8'b00011110;     //219pi/512
   m_sin[220]  =  8'b11001000;     //220pi/512
   m_cos[220]  =  8'b00011110;     //220pi/512
   m_sin[221]  =  8'b11000111;     //221pi/512
   m_cos[221]  =  8'b00011101;     //221pi/512
   m_sin[222]  =  8'b11000111;     //222pi/512
   m_cos[222]  =  8'b00011101;     //222pi/512
   m_sin[223]  =  8'b11000111;     //223pi/512
   m_cos[223]  =  8'b00011101;     //223pi/512
   m_sin[224]  =  8'b11000111;     //224pi/512
   m_cos[224]  =  8'b00011101;     //224pi/512
   m_sin[225]  =  8'b11000111;     //225pi/512
   m_cos[225]  =  8'b00011100;     //225pi/512
   m_sin[226]  =  8'b11000111;     //226pi/512
   m_cos[226]  =  8'b00011100;     //226pi/512
   m_sin[227]  =  8'b11000111;     //227pi/512
   m_cos[227]  =  8'b00011100;     //227pi/512
   m_sin[228]  =  8'b11000110;     //228pi/512
   m_cos[228]  =  8'b00011011;     //228pi/512
   m_sin[229]  =  8'b11000110;     //229pi/512
   m_cos[229]  =  8'b00011011;     //229pi/512
   m_sin[230]  =  8'b11000110;     //230pi/512
   m_cos[230]  =  8'b00011011;     //230pi/512
   m_sin[231]  =  8'b11000110;     //231pi/512
   m_cos[231]  =  8'b00011011;     //231pi/512
   m_sin[232]  =  8'b11000110;     //232pi/512
   m_cos[232]  =  8'b00011010;     //232pi/512
   m_sin[233]  =  8'b11000110;     //233pi/512
   m_cos[233]  =  8'b00011010;     //233pi/512
   m_sin[234]  =  8'b11000110;     //234pi/512
   m_cos[234]  =  8'b00011010;     //234pi/512
   m_sin[235]  =  8'b11000101;     //235pi/512
   m_cos[235]  =  8'b00011001;     //235pi/512
   m_sin[236]  =  8'b11000101;     //236pi/512
   m_cos[236]  =  8'b00011001;     //236pi/512
   m_sin[237]  =  8'b11000101;     //237pi/512
   m_cos[237]  =  8'b00011001;     //237pi/512
   m_sin[238]  =  8'b11000101;     //238pi/512
   m_cos[238]  =  8'b00011001;     //238pi/512
   m_sin[239]  =  8'b11000101;     //239pi/512
   m_cos[239]  =  8'b00011000;     //239pi/512
   m_sin[240]  =  8'b11000101;     //240pi/512
   m_cos[240]  =  8'b00011000;     //240pi/512
   m_sin[241]  =  8'b11000101;     //241pi/512
   m_cos[241]  =  8'b00011000;     //241pi/512
   m_sin[242]  =  8'b11000101;     //242pi/512
   m_cos[242]  =  8'b00010111;     //242pi/512
   m_sin[243]  =  8'b11000101;     //243pi/512
   m_cos[243]  =  8'b00010111;     //243pi/512
   m_sin[244]  =  8'b11000100;     //244pi/512
   m_cos[244]  =  8'b00010111;     //244pi/512
   m_sin[245]  =  8'b11000100;     //245pi/512
   m_cos[245]  =  8'b00010111;     //245pi/512
   m_sin[246]  =  8'b11000100;     //246pi/512
   m_cos[246]  =  8'b00010110;     //246pi/512
   m_sin[247]  =  8'b11000100;     //247pi/512
   m_cos[247]  =  8'b00010110;     //247pi/512
   m_sin[248]  =  8'b11000100;     //248pi/512
   m_cos[248]  =  8'b00010110;     //248pi/512
   m_sin[249]  =  8'b11000100;     //249pi/512
   m_cos[249]  =  8'b00010101;     //249pi/512
   m_sin[250]  =  8'b11000100;     //250pi/512
   m_cos[250]  =  8'b00010101;     //250pi/512
   m_sin[251]  =  8'b11000100;     //251pi/512
   m_cos[251]  =  8'b00010101;     //251pi/512
   m_sin[252]  =  8'b11000100;     //252pi/512
   m_cos[252]  =  8'b00010100;     //252pi/512
   m_sin[253]  =  8'b11000011;     //253pi/512
   m_cos[253]  =  8'b00010100;     //253pi/512
   m_sin[254]  =  8'b11000011;     //254pi/512
   m_cos[254]  =  8'b00010100;     //254pi/512
   m_sin[255]  =  8'b11000011;     //255pi/512
   m_cos[255]  =  8'b00010100;     //255pi/512
   m_sin[256]  =  8'b11000011;     //256pi/512
   m_cos[256]  =  8'b00010011;     //256pi/512
   m_sin[257]  =  8'b11000011;     //257pi/512
   m_cos[257]  =  8'b00010011;     //257pi/512
   m_sin[258]  =  8'b11000011;     //258pi/512
   m_cos[258]  =  8'b00010011;     //258pi/512
   m_sin[259]  =  8'b11000011;     //259pi/512
   m_cos[259]  =  8'b00010010;     //259pi/512
   m_sin[260]  =  8'b11000011;     //260pi/512
   m_cos[260]  =  8'b00010010;     //260pi/512
   m_sin[261]  =  8'b11000011;     //261pi/512
   m_cos[261]  =  8'b00010010;     //261pi/512
   m_sin[262]  =  8'b11000011;     //262pi/512
   m_cos[262]  =  8'b00010001;     //262pi/512
   m_sin[263]  =  8'b11000010;     //263pi/512
   m_cos[263]  =  8'b00010001;     //263pi/512
   m_sin[264]  =  8'b11000010;     //264pi/512
   m_cos[264]  =  8'b00010001;     //264pi/512
   m_sin[265]  =  8'b11000010;     //265pi/512
   m_cos[265]  =  8'b00010001;     //265pi/512
   m_sin[266]  =  8'b11000010;     //266pi/512
   m_cos[266]  =  8'b00010000;     //266pi/512
   m_sin[267]  =  8'b11000010;     //267pi/512
   m_cos[267]  =  8'b00010000;     //267pi/512
   m_sin[268]  =  8'b11000010;     //268pi/512
   m_cos[268]  =  8'b00010000;     //268pi/512
   m_sin[269]  =  8'b11000010;     //269pi/512
   m_cos[269]  =  8'b00001111;     //269pi/512
   m_sin[270]  =  8'b11000010;     //270pi/512
   m_cos[270]  =  8'b00001111;     //270pi/512
   m_sin[271]  =  8'b11000010;     //271pi/512
   m_cos[271]  =  8'b00001111;     //271pi/512
   m_sin[272]  =  8'b11000010;     //272pi/512
   m_cos[272]  =  8'b00001110;     //272pi/512
   m_sin[273]  =  8'b11000010;     //273pi/512
   m_cos[273]  =  8'b00001110;     //273pi/512
   m_sin[274]  =  8'b11000010;     //274pi/512
   m_cos[274]  =  8'b00001110;     //274pi/512
   m_sin[275]  =  8'b11000010;     //275pi/512
   m_cos[275]  =  8'b00001110;     //275pi/512
   m_sin[276]  =  8'b11000001;     //276pi/512
   m_cos[276]  =  8'b00001101;     //276pi/512
   m_sin[277]  =  8'b11000001;     //277pi/512
   m_cos[277]  =  8'b00001101;     //277pi/512
   m_sin[278]  =  8'b11000001;     //278pi/512
   m_cos[278]  =  8'b00001101;     //278pi/512
   m_sin[279]  =  8'b11000001;     //279pi/512
   m_cos[279]  =  8'b00001100;     //279pi/512
   m_sin[280]  =  8'b11000001;     //280pi/512
   m_cos[280]  =  8'b00001100;     //280pi/512
   m_sin[281]  =  8'b11000001;     //281pi/512
   m_cos[281]  =  8'b00001100;     //281pi/512
   m_sin[282]  =  8'b11000001;     //282pi/512
   m_cos[282]  =  8'b00001011;     //282pi/512
   m_sin[283]  =  8'b11000001;     //283pi/512
   m_cos[283]  =  8'b00001011;     //283pi/512
   m_sin[284]  =  8'b11000001;     //284pi/512
   m_cos[284]  =  8'b00001011;     //284pi/512
   m_sin[285]  =  8'b11000001;     //285pi/512
   m_cos[285]  =  8'b00001010;     //285pi/512
   m_sin[286]  =  8'b11000001;     //286pi/512
   m_cos[286]  =  8'b00001010;     //286pi/512
   m_sin[287]  =  8'b11000001;     //287pi/512
   m_cos[287]  =  8'b00001010;     //287pi/512
   m_sin[288]  =  8'b11000001;     //288pi/512
   m_cos[288]  =  8'b00001010;     //288pi/512
   m_sin[289]  =  8'b11000001;     //289pi/512
   m_cos[289]  =  8'b00001001;     //289pi/512
   m_sin[290]  =  8'b11000001;     //290pi/512
   m_cos[290]  =  8'b00001001;     //290pi/512
   m_sin[291]  =  8'b11000001;     //291pi/512
   m_cos[291]  =  8'b00001001;     //291pi/512
   m_sin[292]  =  8'b11000001;     //292pi/512
   m_cos[292]  =  8'b00001000;     //292pi/512
   m_sin[293]  =  8'b11000001;     //293pi/512
   m_cos[293]  =  8'b00001000;     //293pi/512
   m_sin[294]  =  8'b11000001;     //294pi/512
   m_cos[294]  =  8'b00001000;     //294pi/512
   m_sin[295]  =  8'b11000000;     //295pi/512
   m_cos[295]  =  8'b00000111;     //295pi/512
   m_sin[296]  =  8'b11000000;     //296pi/512
   m_cos[296]  =  8'b00000111;     //296pi/512
   m_sin[297]  =  8'b11000000;     //297pi/512
   m_cos[297]  =  8'b00000111;     //297pi/512
   m_sin[298]  =  8'b11000000;     //298pi/512
   m_cos[298]  =  8'b00000110;     //298pi/512
   m_sin[299]  =  8'b11000000;     //299pi/512
   m_cos[299]  =  8'b00000110;     //299pi/512
   m_sin[300]  =  8'b11000000;     //300pi/512
   m_cos[300]  =  8'b00000110;     //300pi/512
   m_sin[301]  =  8'b11000000;     //301pi/512
   m_cos[301]  =  8'b00000101;     //301pi/512
   m_sin[302]  =  8'b11000000;     //302pi/512
   m_cos[302]  =  8'b00000101;     //302pi/512
   m_sin[303]  =  8'b11000000;     //303pi/512
   m_cos[303]  =  8'b00000101;     //303pi/512
   m_sin[304]  =  8'b11000000;     //304pi/512
   m_cos[304]  =  8'b00000101;     //304pi/512
   m_sin[305]  =  8'b11000000;     //305pi/512
   m_cos[305]  =  8'b00000100;     //305pi/512
   m_sin[306]  =  8'b11000000;     //306pi/512
   m_cos[306]  =  8'b00000100;     //306pi/512
   m_sin[307]  =  8'b11000000;     //307pi/512
   m_cos[307]  =  8'b00000100;     //307pi/512
   m_sin[308]  =  8'b11000000;     //308pi/512
   m_cos[308]  =  8'b00000011;     //308pi/512
   m_sin[309]  =  8'b11000000;     //309pi/512
   m_cos[309]  =  8'b00000011;     //309pi/512
   m_sin[310]  =  8'b11000000;     //310pi/512
   m_cos[310]  =  8'b00000011;     //310pi/512
   m_sin[311]  =  8'b11000000;     //311pi/512
   m_cos[311]  =  8'b00000010;     //311pi/512
   m_sin[312]  =  8'b11000000;     //312pi/512
   m_cos[312]  =  8'b00000010;     //312pi/512
   m_sin[313]  =  8'b11000000;     //313pi/512
   m_cos[313]  =  8'b00000010;     //313pi/512
   m_sin[314]  =  8'b11000000;     //314pi/512
   m_cos[314]  =  8'b00000001;     //314pi/512
   m_sin[315]  =  8'b11000000;     //315pi/512
   m_cos[315]  =  8'b00000001;     //315pi/512
   m_sin[316]  =  8'b11000000;     //316pi/512
   m_cos[316]  =  8'b00000001;     //316pi/512
   m_sin[317]  =  8'b11000000;     //317pi/512
   m_cos[317]  =  8'b00000000;     //317pi/512
   m_sin[318]  =  8'b11000000;     //318pi/512
   m_cos[318]  =  8'b00000000;     //318pi/512
   m_sin[319]  =  8'b11000000;     //319pi/512
   m_cos[319]  =  8'b00000000;     //319pi/512
   m_sin[320]  =  8'b11000000;     //320pi/512
   m_cos[320]  =  8'b00000000;     //320pi/512
   m_sin[321]  =  8'b11000000;     //321pi/512
   m_cos[321]  =  8'b00000000;     //321pi/512
   m_sin[322]  =  8'b11000000;     //322pi/512
   m_cos[322]  =  8'b11111111;     //322pi/512
   m_sin[323]  =  8'b11000000;     //323pi/512
   m_cos[323]  =  8'b11111111;     //323pi/512
   m_sin[324]  =  8'b11000000;     //324pi/512
   m_cos[324]  =  8'b11111111;     //324pi/512
   m_sin[325]  =  8'b11000000;     //325pi/512
   m_cos[325]  =  8'b11111110;     //325pi/512
   m_sin[326]  =  8'b11000000;     //326pi/512
   m_cos[326]  =  8'b11111110;     //326pi/512
   m_sin[327]  =  8'b11000000;     //327pi/512
   m_cos[327]  =  8'b11111110;     //327pi/512
   m_sin[328]  =  8'b11000000;     //328pi/512
   m_cos[328]  =  8'b11111101;     //328pi/512
   m_sin[329]  =  8'b11000000;     //329pi/512
   m_cos[329]  =  8'b11111101;     //329pi/512
   m_sin[330]  =  8'b11000000;     //330pi/512
   m_cos[330]  =  8'b11111101;     //330pi/512
   m_sin[331]  =  8'b11000000;     //331pi/512
   m_cos[331]  =  8'b11111101;     //331pi/512
   m_sin[332]  =  8'b11000000;     //332pi/512
   m_cos[332]  =  8'b11111100;     //332pi/512
   m_sin[333]  =  8'b11000000;     //333pi/512
   m_cos[333]  =  8'b11111100;     //333pi/512
   m_sin[334]  =  8'b11000000;     //334pi/512
   m_cos[334]  =  8'b11111100;     //334pi/512
   m_sin[335]  =  8'b11000000;     //335pi/512
   m_cos[335]  =  8'b11111011;     //335pi/512
   m_sin[336]  =  8'b11000000;     //336pi/512
   m_cos[336]  =  8'b11111011;     //336pi/512
   m_sin[337]  =  8'b11000000;     //337pi/512
   m_cos[337]  =  8'b11111011;     //337pi/512
   m_sin[338]  =  8'b11000000;     //338pi/512
   m_cos[338]  =  8'b11111010;     //338pi/512
   m_sin[339]  =  8'b11000000;     //339pi/512
   m_cos[339]  =  8'b11111010;     //339pi/512
   m_sin[340]  =  8'b11000000;     //340pi/512
   m_cos[340]  =  8'b11111010;     //340pi/512
   m_sin[341]  =  8'b11000000;     //341pi/512
   m_cos[341]  =  8'b11111001;     //341pi/512
   m_sin[342]  =  8'b11000000;     //342pi/512
   m_cos[342]  =  8'b11111001;     //342pi/512
   m_sin[343]  =  8'b11000000;     //343pi/512
   m_cos[343]  =  8'b11111001;     //343pi/512
   m_sin[344]  =  8'b11000000;     //344pi/512
   m_cos[344]  =  8'b11111000;     //344pi/512
   m_sin[345]  =  8'b11000000;     //345pi/512
   m_cos[345]  =  8'b11111000;     //345pi/512
   m_sin[346]  =  8'b11000001;     //346pi/512
   m_cos[346]  =  8'b11111000;     //346pi/512
   m_sin[347]  =  8'b11000001;     //347pi/512
   m_cos[347]  =  8'b11111000;     //347pi/512
   m_sin[348]  =  8'b11000001;     //348pi/512
   m_cos[348]  =  8'b11110111;     //348pi/512
   m_sin[349]  =  8'b11000001;     //349pi/512
   m_cos[349]  =  8'b11110111;     //349pi/512
   m_sin[350]  =  8'b11000001;     //350pi/512
   m_cos[350]  =  8'b11110111;     //350pi/512
   m_sin[351]  =  8'b11000001;     //351pi/512
   m_cos[351]  =  8'b11110110;     //351pi/512
   m_sin[352]  =  8'b11000001;     //352pi/512
   m_cos[352]  =  8'b11110110;     //352pi/512
   m_sin[353]  =  8'b11000001;     //353pi/512
   m_cos[353]  =  8'b11110110;     //353pi/512
   m_sin[354]  =  8'b11000001;     //354pi/512
   m_cos[354]  =  8'b11110101;     //354pi/512
   m_sin[355]  =  8'b11000001;     //355pi/512
   m_cos[355]  =  8'b11110101;     //355pi/512
   m_sin[356]  =  8'b11000001;     //356pi/512
   m_cos[356]  =  8'b11110101;     //356pi/512
   m_sin[357]  =  8'b11000001;     //357pi/512
   m_cos[357]  =  8'b11110100;     //357pi/512
   m_sin[358]  =  8'b11000001;     //358pi/512
   m_cos[358]  =  8'b11110100;     //358pi/512
   m_sin[359]  =  8'b11000001;     //359pi/512
   m_cos[359]  =  8'b11110100;     //359pi/512
   m_sin[360]  =  8'b11000001;     //360pi/512
   m_cos[360]  =  8'b11110100;     //360pi/512
   m_sin[361]  =  8'b11000001;     //361pi/512
   m_cos[361]  =  8'b11110011;     //361pi/512
   m_sin[362]  =  8'b11000001;     //362pi/512
   m_cos[362]  =  8'b11110011;     //362pi/512
   m_sin[363]  =  8'b11000001;     //363pi/512
   m_cos[363]  =  8'b11110011;     //363pi/512
   m_sin[364]  =  8'b11000001;     //364pi/512
   m_cos[364]  =  8'b11110010;     //364pi/512
   m_sin[365]  =  8'b11000010;     //365pi/512
   m_cos[365]  =  8'b11110010;     //365pi/512
   m_sin[366]  =  8'b11000010;     //366pi/512
   m_cos[366]  =  8'b11110010;     //366pi/512
   m_sin[367]  =  8'b11000010;     //367pi/512
   m_cos[367]  =  8'b11110001;     //367pi/512
   m_sin[368]  =  8'b11000010;     //368pi/512
   m_cos[368]  =  8'b11110001;     //368pi/512
   m_sin[369]  =  8'b11000010;     //369pi/512
   m_cos[369]  =  8'b11110001;     //369pi/512
   m_sin[370]  =  8'b11000010;     //370pi/512
   m_cos[370]  =  8'b11110000;     //370pi/512
   m_sin[371]  =  8'b11000010;     //371pi/512
   m_cos[371]  =  8'b11110000;     //371pi/512
   m_sin[372]  =  8'b11000010;     //372pi/512
   m_cos[372]  =  8'b11110000;     //372pi/512
   m_sin[373]  =  8'b11000010;     //373pi/512
   m_cos[373]  =  8'b11110000;     //373pi/512
   m_sin[374]  =  8'b11000010;     //374pi/512
   m_cos[374]  =  8'b11101111;     //374pi/512
   m_sin[375]  =  8'b11000010;     //375pi/512
   m_cos[375]  =  8'b11101111;     //375pi/512
   m_sin[376]  =  8'b11000010;     //376pi/512
   m_cos[376]  =  8'b11101111;     //376pi/512
   m_sin[377]  =  8'b11000010;     //377pi/512
   m_cos[377]  =  8'b11101110;     //377pi/512
   m_sin[378]  =  8'b11000011;     //378pi/512
   m_cos[378]  =  8'b11101110;     //378pi/512
   m_sin[379]  =  8'b11000011;     //379pi/512
   m_cos[379]  =  8'b11101110;     //379pi/512
   m_sin[380]  =  8'b11000011;     //380pi/512
   m_cos[380]  =  8'b11101101;     //380pi/512
   m_sin[381]  =  8'b11000011;     //381pi/512
   m_cos[381]  =  8'b11101101;     //381pi/512
   m_sin[382]  =  8'b11000011;     //382pi/512
   m_cos[382]  =  8'b11101101;     //382pi/512
   m_sin[383]  =  8'b11000011;     //383pi/512
   m_cos[383]  =  8'b11101101;     //383pi/512
   m_sin[384]  =  8'b11000011;     //384pi/512
   m_cos[384]  =  8'b11101100;     //384pi/512
   m_sin[385]  =  8'b11000011;     //385pi/512
   m_cos[385]  =  8'b11101100;     //385pi/512
   m_sin[386]  =  8'b11000011;     //386pi/512
   m_cos[386]  =  8'b11101100;     //386pi/512
   m_sin[387]  =  8'b11000011;     //387pi/512
   m_cos[387]  =  8'b11101011;     //387pi/512
   m_sin[388]  =  8'b11000100;     //388pi/512
   m_cos[388]  =  8'b11101011;     //388pi/512
   m_sin[389]  =  8'b11000100;     //389pi/512
   m_cos[389]  =  8'b11101011;     //389pi/512
   m_sin[390]  =  8'b11000100;     //390pi/512
   m_cos[390]  =  8'b11101010;     //390pi/512
   m_sin[391]  =  8'b11000100;     //391pi/512
   m_cos[391]  =  8'b11101010;     //391pi/512
   m_sin[392]  =  8'b11000100;     //392pi/512
   m_cos[392]  =  8'b11101010;     //392pi/512
   m_sin[393]  =  8'b11000100;     //393pi/512
   m_cos[393]  =  8'b11101010;     //393pi/512
   m_sin[394]  =  8'b11000100;     //394pi/512
   m_cos[394]  =  8'b11101001;     //394pi/512
   m_sin[395]  =  8'b11000100;     //395pi/512
   m_cos[395]  =  8'b11101001;     //395pi/512
   m_sin[396]  =  8'b11000100;     //396pi/512
   m_cos[396]  =  8'b11101001;     //396pi/512
   m_sin[397]  =  8'b11000101;     //397pi/512
   m_cos[397]  =  8'b11101000;     //397pi/512
   m_sin[398]  =  8'b11000101;     //398pi/512
   m_cos[398]  =  8'b11101000;     //398pi/512
   m_sin[399]  =  8'b11000101;     //399pi/512
   m_cos[399]  =  8'b11101000;     //399pi/512
   m_sin[400]  =  8'b11000101;     //400pi/512
   m_cos[400]  =  8'b11101000;     //400pi/512
   m_sin[401]  =  8'b11000101;     //401pi/512
   m_cos[401]  =  8'b11100111;     //401pi/512
   m_sin[402]  =  8'b11000101;     //402pi/512
   m_cos[402]  =  8'b11100111;     //402pi/512
   m_sin[403]  =  8'b11000101;     //403pi/512
   m_cos[403]  =  8'b11100111;     //403pi/512
   m_sin[404]  =  8'b11000101;     //404pi/512
   m_cos[404]  =  8'b11100110;     //404pi/512
   m_sin[405]  =  8'b11000101;     //405pi/512
   m_cos[405]  =  8'b11100110;     //405pi/512
   m_sin[406]  =  8'b11000110;     //406pi/512
   m_cos[406]  =  8'b11100110;     //406pi/512
   m_sin[407]  =  8'b11000110;     //407pi/512
   m_cos[407]  =  8'b11100101;     //407pi/512
   m_sin[408]  =  8'b11000110;     //408pi/512
   m_cos[408]  =  8'b11100101;     //408pi/512
   m_sin[409]  =  8'b11000110;     //409pi/512
   m_cos[409]  =  8'b11100101;     //409pi/512
   m_sin[410]  =  8'b11000110;     //410pi/512
   m_cos[410]  =  8'b11100101;     //410pi/512
   m_sin[411]  =  8'b11000110;     //411pi/512
   m_cos[411]  =  8'b11100100;     //411pi/512
   m_sin[412]  =  8'b11000110;     //412pi/512
   m_cos[412]  =  8'b11100100;     //412pi/512
   m_sin[413]  =  8'b11000111;     //413pi/512
   m_cos[413]  =  8'b11100100;     //413pi/512
   m_sin[414]  =  8'b11000111;     //414pi/512
   m_cos[414]  =  8'b11100100;     //414pi/512
   m_sin[415]  =  8'b11000111;     //415pi/512
   m_cos[415]  =  8'b11100011;     //415pi/512
   m_sin[416]  =  8'b11000111;     //416pi/512
   m_cos[416]  =  8'b11100011;     //416pi/512
   m_sin[417]  =  8'b11000111;     //417pi/512
   m_cos[417]  =  8'b11100011;     //417pi/512
   m_sin[418]  =  8'b11000111;     //418pi/512
   m_cos[418]  =  8'b11100010;     //418pi/512
   m_sin[419]  =  8'b11000111;     //419pi/512
   m_cos[419]  =  8'b11100010;     //419pi/512
   m_sin[420]  =  8'b11001000;     //420pi/512
   m_cos[420]  =  8'b11100010;     //420pi/512
   m_sin[421]  =  8'b11001000;     //421pi/512
   m_cos[421]  =  8'b11100010;     //421pi/512
   m_sin[422]  =  8'b11001000;     //422pi/512
   m_cos[422]  =  8'b11100001;     //422pi/512
   m_sin[423]  =  8'b11001000;     //423pi/512
   m_cos[423]  =  8'b11100001;     //423pi/512
   m_sin[424]  =  8'b11001000;     //424pi/512
   m_cos[424]  =  8'b11100001;     //424pi/512
   m_sin[425]  =  8'b11001000;     //425pi/512
   m_cos[425]  =  8'b11100000;     //425pi/512
   m_sin[426]  =  8'b11001000;     //426pi/512
   m_cos[426]  =  8'b11100000;     //426pi/512
   m_sin[427]  =  8'b11001001;     //427pi/512
   m_cos[427]  =  8'b11100000;     //427pi/512
   m_sin[428]  =  8'b11001001;     //428pi/512
   m_cos[428]  =  8'b11100000;     //428pi/512
   m_sin[429]  =  8'b11001001;     //429pi/512
   m_cos[429]  =  8'b11011111;     //429pi/512
   m_sin[430]  =  8'b11001001;     //430pi/512
   m_cos[430]  =  8'b11011111;     //430pi/512
   m_sin[431]  =  8'b11001001;     //431pi/512
   m_cos[431]  =  8'b11011111;     //431pi/512
   m_sin[432]  =  8'b11001001;     //432pi/512
   m_cos[432]  =  8'b11011111;     //432pi/512
   m_sin[433]  =  8'b11001010;     //433pi/512
   m_cos[433]  =  8'b11011110;     //433pi/512
   m_sin[434]  =  8'b11001010;     //434pi/512
   m_cos[434]  =  8'b11011110;     //434pi/512
   m_sin[435]  =  8'b11001010;     //435pi/512
   m_cos[435]  =  8'b11011110;     //435pi/512
   m_sin[436]  =  8'b11001010;     //436pi/512
   m_cos[436]  =  8'b11011101;     //436pi/512
   m_sin[437]  =  8'b11001010;     //437pi/512
   m_cos[437]  =  8'b11011101;     //437pi/512
   m_sin[438]  =  8'b11001010;     //438pi/512
   m_cos[438]  =  8'b11011101;     //438pi/512
   m_sin[439]  =  8'b11001011;     //439pi/512
   m_cos[439]  =  8'b11011101;     //439pi/512
   m_sin[440]  =  8'b11001011;     //440pi/512
   m_cos[440]  =  8'b11011100;     //440pi/512
   m_sin[441]  =  8'b11001011;     //441pi/512
   m_cos[441]  =  8'b11011100;     //441pi/512
   m_sin[442]  =  8'b11001011;     //442pi/512
   m_cos[442]  =  8'b11011100;     //442pi/512
   m_sin[443]  =  8'b11001011;     //443pi/512
   m_cos[443]  =  8'b11011100;     //443pi/512
   m_sin[444]  =  8'b11001011;     //444pi/512
   m_cos[444]  =  8'b11011011;     //444pi/512
   m_sin[445]  =  8'b11001100;     //445pi/512
   m_cos[445]  =  8'b11011011;     //445pi/512
   m_sin[446]  =  8'b11001100;     //446pi/512
   m_cos[446]  =  8'b11011011;     //446pi/512
   m_sin[447]  =  8'b11001100;     //447pi/512
   m_cos[447]  =  8'b11011011;     //447pi/512
   m_sin[448]  =  8'b11001100;     //448pi/512
   m_cos[448]  =  8'b11011010;     //448pi/512
   m_sin[449]  =  8'b11001100;     //449pi/512
   m_cos[449]  =  8'b11011010;     //449pi/512
   m_sin[450]  =  8'b11001101;     //450pi/512
   m_cos[450]  =  8'b11011010;     //450pi/512
   m_sin[451]  =  8'b11001101;     //451pi/512
   m_cos[451]  =  8'b11011010;     //451pi/512
   m_sin[452]  =  8'b11001101;     //452pi/512
   m_cos[452]  =  8'b11011001;     //452pi/512
   m_sin[453]  =  8'b11001101;     //453pi/512
   m_cos[453]  =  8'b11011001;     //453pi/512
   m_sin[454]  =  8'b11001101;     //454pi/512
   m_cos[454]  =  8'b11011001;     //454pi/512
   m_sin[455]  =  8'b11001110;     //455pi/512
   m_cos[455]  =  8'b11011001;     //455pi/512
   m_sin[456]  =  8'b11001110;     //456pi/512
   m_cos[456]  =  8'b11011000;     //456pi/512
   m_sin[457]  =  8'b11001110;     //457pi/512
   m_cos[457]  =  8'b11011000;     //457pi/512
   m_sin[458]  =  8'b11001110;     //458pi/512
   m_cos[458]  =  8'b11011000;     //458pi/512
   m_sin[459]  =  8'b11001110;     //459pi/512
   m_cos[459]  =  8'b11011000;     //459pi/512
   m_sin[460]  =  8'b11001111;     //460pi/512
   m_cos[460]  =  8'b11010111;     //460pi/512
   m_sin[461]  =  8'b11001111;     //461pi/512
   m_cos[461]  =  8'b11010111;     //461pi/512
   m_sin[462]  =  8'b11001111;     //462pi/512
   m_cos[462]  =  8'b11010111;     //462pi/512
   m_sin[463]  =  8'b11001111;     //463pi/512
   m_cos[463]  =  8'b11010111;     //463pi/512
   m_sin[464]  =  8'b11001111;     //464pi/512
   m_cos[464]  =  8'b11010110;     //464pi/512
   m_sin[465]  =  8'b11010000;     //465pi/512
   m_cos[465]  =  8'b11010110;     //465pi/512
   m_sin[466]  =  8'b11010000;     //466pi/512
   m_cos[466]  =  8'b11010110;     //466pi/512
   m_sin[467]  =  8'b11010000;     //467pi/512
   m_cos[467]  =  8'b11010110;     //467pi/512
   m_sin[468]  =  8'b11010000;     //468pi/512
   m_cos[468]  =  8'b11010101;     //468pi/512
   m_sin[469]  =  8'b11010000;     //469pi/512
   m_cos[469]  =  8'b11010101;     //469pi/512
   m_sin[470]  =  8'b11010001;     //470pi/512
   m_cos[470]  =  8'b11010101;     //470pi/512
   m_sin[471]  =  8'b11010001;     //471pi/512
   m_cos[471]  =  8'b11010101;     //471pi/512
   m_sin[472]  =  8'b11010001;     //472pi/512
   m_cos[472]  =  8'b11010101;     //472pi/512
   m_sin[473]  =  8'b11010001;     //473pi/512
   m_cos[473]  =  8'b11010100;     //473pi/512
   m_sin[474]  =  8'b11010001;     //474pi/512
   m_cos[474]  =  8'b11010100;     //474pi/512
   m_sin[475]  =  8'b11010010;     //475pi/512
   m_cos[475]  =  8'b11010100;     //475pi/512
   m_sin[476]  =  8'b11010010;     //476pi/512
   m_cos[476]  =  8'b11010100;     //476pi/512
   m_sin[477]  =  8'b11010010;     //477pi/512
   m_cos[477]  =  8'b11010011;     //477pi/512
   m_sin[478]  =  8'b11010010;     //478pi/512
   m_cos[478]  =  8'b11010011;     //478pi/512
   m_sin[479]  =  8'b11010011;     //479pi/512
   m_cos[479]  =  8'b11010011;     //479pi/512
   m_sin[480]  =  8'b11010011;     //480pi/512
   m_cos[480]  =  8'b11010011;     //480pi/512
   m_sin[481]  =  8'b11010011;     //481pi/512
   m_cos[481]  =  8'b11010011;     //481pi/512
   m_sin[482]  =  8'b11010011;     //482pi/512
   m_cos[482]  =  8'b11010010;     //482pi/512
   m_sin[483]  =  8'b11010011;     //483pi/512
   m_cos[483]  =  8'b11010010;     //483pi/512
   m_sin[484]  =  8'b11010100;     //484pi/512
   m_cos[484]  =  8'b11010010;     //484pi/512
   m_sin[485]  =  8'b11010100;     //485pi/512
   m_cos[485]  =  8'b11010010;     //485pi/512
   m_sin[486]  =  8'b11010100;     //486pi/512
   m_cos[486]  =  8'b11010001;     //486pi/512
   m_sin[487]  =  8'b11010100;     //487pi/512
   m_cos[487]  =  8'b11010001;     //487pi/512
   m_sin[488]  =  8'b11010101;     //488pi/512
   m_cos[488]  =  8'b11010001;     //488pi/512
   m_sin[489]  =  8'b11010101;     //489pi/512
   m_cos[489]  =  8'b11010001;     //489pi/512
   m_sin[490]  =  8'b11010101;     //490pi/512
   m_cos[490]  =  8'b11010001;     //490pi/512
   m_sin[491]  =  8'b11010101;     //491pi/512
   m_cos[491]  =  8'b11010000;     //491pi/512
   m_sin[492]  =  8'b11010101;     //492pi/512
   m_cos[492]  =  8'b11010000;     //492pi/512
   m_sin[493]  =  8'b11010110;     //493pi/512
   m_cos[493]  =  8'b11010000;     //493pi/512
   m_sin[494]  =  8'b11010110;     //494pi/512
   m_cos[494]  =  8'b11010000;     //494pi/512
   m_sin[495]  =  8'b11010110;     //495pi/512
   m_cos[495]  =  8'b11010000;     //495pi/512
   m_sin[496]  =  8'b11010110;     //496pi/512
   m_cos[496]  =  8'b11001111;     //496pi/512
   m_sin[497]  =  8'b11010111;     //497pi/512
   m_cos[497]  =  8'b11001111;     //497pi/512
   m_sin[498]  =  8'b11010111;     //498pi/512
   m_cos[498]  =  8'b11001111;     //498pi/512
   m_sin[499]  =  8'b11010111;     //499pi/512
   m_cos[499]  =  8'b11001111;     //499pi/512
   m_sin[500]  =  8'b11010111;     //500pi/512
   m_cos[500]  =  8'b11001111;     //500pi/512
   m_sin[501]  =  8'b11011000;     //501pi/512
   m_cos[501]  =  8'b11001110;     //501pi/512
   m_sin[502]  =  8'b11011000;     //502pi/512
   m_cos[502]  =  8'b11001110;     //502pi/512
   m_sin[503]  =  8'b11011000;     //503pi/512
   m_cos[503]  =  8'b11001110;     //503pi/512
   m_sin[504]  =  8'b11011000;     //504pi/512
   m_cos[504]  =  8'b11001110;     //504pi/512
   m_sin[505]  =  8'b11011001;     //505pi/512
   m_cos[505]  =  8'b11001110;     //505pi/512
   m_sin[506]  =  8'b11011001;     //506pi/512
   m_cos[506]  =  8'b11001101;     //506pi/512
   m_sin[507]  =  8'b11011001;     //507pi/512
   m_cos[507]  =  8'b11001101;     //507pi/512
   m_sin[508]  =  8'b11011001;     //508pi/512
   m_cos[508]  =  8'b11001101;     //508pi/512
   m_sin[509]  =  8'b11011010;     //509pi/512
   m_cos[509]  =  8'b11001101;     //509pi/512
   m_sin[510]  =  8'b11011010;     //510pi/512
   m_cos[510]  =  8'b11001101;     //510pi/512
   m_sin[511]  =  8'b11011010;     //511pi/512
   m_cos[511]  =  8'b11001100;     //511pi/512
end
endmodule