module  M_TWIDLE_7_bit #(parameter SIZE =10) (
    input            en_modify, 
    input   [10:0]   rd_ptr_angle,

    output  signed [6:0]   cos_data,
    output  signed [6:0]   sin_data
 );


wire signed [6:0]  cos  [511:0];
wire signed [6:0]  sin  [511:0];

wire signed [6:0]  cos2  [511:0];
wire signed [6:0]  sin2  [511:0];

assign cos_data =   en_modify? cos2 [rd_ptr_angle] : cos [rd_ptr_angle];
assign sin_data =   en_modify? sin2 [rd_ptr_angle] : sin [rd_ptr_angle];

  assign sin[0]  =  7'b0000000;     //0pi/512
  assign cos[0]  =  7'b0100000;     //0pi/512
  assign sin[1]  =  7'b0000000;     //1pi/512
  assign cos[1]  =  7'b0011111;     //1pi/512
  assign sin[2]  =  7'b0000000;     //2pi/512
  assign cos[2]  =  7'b0011111;     //2pi/512
  assign sin[3]  =  7'b1111111;     //3pi/512
  assign cos[3]  =  7'b0011111;     //3pi/512
  assign sin[4]  =  7'b1111111;     //4pi/512
  assign cos[4]  =  7'b0011111;     //4pi/512
  assign sin[5]  =  7'b1111111;     //5pi/512
  assign cos[5]  =  7'b0011111;     //5pi/512
  assign sin[6]  =  7'b1111111;     //6pi/512
  assign cos[6]  =  7'b0011111;     //6pi/512
  assign sin[7]  =  7'b1111111;     //7pi/512
  assign cos[7]  =  7'b0011111;     //7pi/512
  assign sin[8]  =  7'b1111110;     //8pi/512
  assign cos[8]  =  7'b0011111;     //8pi/512
  assign sin[9]  =  7'b1111110;     //9pi/512
  assign cos[9]  =  7'b0011111;     //9pi/512
  assign sin[10]  =  7'b1111110;     //10pi/512
  assign cos[10]  =  7'b0011111;     //10pi/512
  assign sin[11]  =  7'b1111110;     //11pi/512
  assign cos[11]  =  7'b0011111;     //11pi/512
  assign sin[12]  =  7'b1111110;     //12pi/512
  assign cos[12]  =  7'b0011111;     //12pi/512
  assign sin[13]  =  7'b1111101;     //13pi/512
  assign cos[13]  =  7'b0011111;     //13pi/512
  assign sin[14]  =  7'b1111101;     //14pi/512
  assign cos[14]  =  7'b0011111;     //14pi/512
  assign sin[15]  =  7'b1111101;     //15pi/512
  assign cos[15]  =  7'b0011111;     //15pi/512
  assign sin[16]  =  7'b1111101;     //16pi/512
  assign cos[16]  =  7'b0011111;     //16pi/512
  assign sin[17]  =  7'b1111101;     //17pi/512
  assign cos[17]  =  7'b0011111;     //17pi/512
  assign sin[18]  =  7'b1111100;     //18pi/512
  assign cos[18]  =  7'b0011111;     //18pi/512
  assign sin[19]  =  7'b1111100;     //19pi/512
  assign cos[19]  =  7'b0011111;     //19pi/512
  assign sin[20]  =  7'b1111100;     //20pi/512
  assign cos[20]  =  7'b0011111;     //20pi/512
  assign sin[21]  =  7'b1111100;     //21pi/512
  assign cos[21]  =  7'b0011111;     //21pi/512
  assign sin[22]  =  7'b1111100;     //22pi/512
  assign cos[22]  =  7'b0011111;     //22pi/512
  assign sin[23]  =  7'b1111011;     //23pi/512
  assign cos[23]  =  7'b0011111;     //23pi/512
  assign sin[24]  =  7'b1111011;     //24pi/512
  assign cos[24]  =  7'b0011111;     //24pi/512
  assign sin[25]  =  7'b1111011;     //25pi/512
  assign cos[25]  =  7'b0011111;     //25pi/512
  assign sin[26]  =  7'b1111011;     //26pi/512
  assign cos[26]  =  7'b0011111;     //26pi/512
  assign sin[27]  =  7'b1111011;     //27pi/512
  assign cos[27]  =  7'b0011111;     //27pi/512
  assign sin[28]  =  7'b1111011;     //28pi/512
  assign cos[28]  =  7'b0011111;     //28pi/512
  assign sin[29]  =  7'b1111010;     //29pi/512
  assign cos[29]  =  7'b0011111;     //29pi/512
  assign sin[30]  =  7'b1111010;     //30pi/512
  assign cos[30]  =  7'b0011111;     //30pi/512
  assign sin[31]  =  7'b1111010;     //31pi/512
  assign cos[31]  =  7'b0011111;     //31pi/512
  assign sin[32]  =  7'b1111010;     //32pi/512
  assign cos[32]  =  7'b0011111;     //32pi/512
  assign sin[33]  =  7'b1111010;     //33pi/512
  assign cos[33]  =  7'b0011111;     //33pi/512
  assign sin[34]  =  7'b1111001;     //34pi/512
  assign cos[34]  =  7'b0011111;     //34pi/512
  assign sin[35]  =  7'b1111001;     //35pi/512
  assign cos[35]  =  7'b0011111;     //35pi/512
  assign sin[36]  =  7'b1111001;     //36pi/512
  assign cos[36]  =  7'b0011111;     //36pi/512
  assign sin[37]  =  7'b1111001;     //37pi/512
  assign cos[37]  =  7'b0011111;     //37pi/512
  assign sin[38]  =  7'b1111001;     //38pi/512
  assign cos[38]  =  7'b0011111;     //38pi/512
  assign sin[39]  =  7'b1111000;     //39pi/512
  assign cos[39]  =  7'b0011111;     //39pi/512
  assign sin[40]  =  7'b1111000;     //40pi/512
  assign cos[40]  =  7'b0011111;     //40pi/512
  assign sin[41]  =  7'b1111000;     //41pi/512
  assign cos[41]  =  7'b0011110;     //41pi/512
  assign sin[42]  =  7'b1111000;     //42pi/512
  assign cos[42]  =  7'b0011110;     //42pi/512
  assign sin[43]  =  7'b1111000;     //43pi/512
  assign cos[43]  =  7'b0011110;     //43pi/512
  assign sin[44]  =  7'b1110111;     //44pi/512
  assign cos[44]  =  7'b0011110;     //44pi/512
  assign sin[45]  =  7'b1110111;     //45pi/512
  assign cos[45]  =  7'b0011110;     //45pi/512
  assign sin[46]  =  7'b1110111;     //46pi/512
  assign cos[46]  =  7'b0011110;     //46pi/512
  assign sin[47]  =  7'b1110111;     //47pi/512
  assign cos[47]  =  7'b0011110;     //47pi/512
  assign sin[48]  =  7'b1110111;     //48pi/512
  assign cos[48]  =  7'b0011110;     //48pi/512
  assign sin[49]  =  7'b1110111;     //49pi/512
  assign cos[49]  =  7'b0011110;     //49pi/512
  assign sin[50]  =  7'b1110110;     //50pi/512
  assign cos[50]  =  7'b0011110;     //50pi/512
  assign sin[51]  =  7'b1110110;     //51pi/512
  assign cos[51]  =  7'b0011110;     //51pi/512
  assign sin[52]  =  7'b1110110;     //52pi/512
  assign cos[52]  =  7'b0011110;     //52pi/512
  assign sin[53]  =  7'b1110110;     //53pi/512
  assign cos[53]  =  7'b0011110;     //53pi/512
  assign sin[54]  =  7'b1110110;     //54pi/512
  assign cos[54]  =  7'b0011110;     //54pi/512
  assign sin[55]  =  7'b1110101;     //55pi/512
  assign cos[55]  =  7'b0011110;     //55pi/512
  assign sin[56]  =  7'b1110101;     //56pi/512
  assign cos[56]  =  7'b0011110;     //56pi/512
  assign sin[57]  =  7'b1110101;     //57pi/512
  assign cos[57]  =  7'b0011110;     //57pi/512
  assign sin[58]  =  7'b1110101;     //58pi/512
  assign cos[58]  =  7'b0011101;     //58pi/512
  assign sin[59]  =  7'b1110101;     //59pi/512
  assign cos[59]  =  7'b0011101;     //59pi/512
  assign sin[60]  =  7'b1110100;     //60pi/512
  assign cos[60]  =  7'b0011101;     //60pi/512
  assign sin[61]  =  7'b1110100;     //61pi/512
  assign cos[61]  =  7'b0011101;     //61pi/512
  assign sin[62]  =  7'b1110100;     //62pi/512
  assign cos[62]  =  7'b0011101;     //62pi/512
  assign sin[63]  =  7'b1110100;     //63pi/512
  assign cos[63]  =  7'b0011101;     //63pi/512
  assign sin[64]  =  7'b1110100;     //64pi/512
  assign cos[64]  =  7'b0011101;     //64pi/512
  assign sin[65]  =  7'b1110100;     //65pi/512
  assign cos[65]  =  7'b0011101;     //65pi/512
  assign sin[66]  =  7'b1110011;     //66pi/512
  assign cos[66]  =  7'b0011101;     //66pi/512
  assign sin[67]  =  7'b1110011;     //67pi/512
  assign cos[67]  =  7'b0011101;     //67pi/512
  assign sin[68]  =  7'b1110011;     //68pi/512
  assign cos[68]  =  7'b0011101;     //68pi/512
  assign sin[69]  =  7'b1110011;     //69pi/512
  assign cos[69]  =  7'b0011101;     //69pi/512
  assign sin[70]  =  7'b1110011;     //70pi/512
  assign cos[70]  =  7'b0011101;     //70pi/512
  assign sin[71]  =  7'b1110010;     //71pi/512
  assign cos[71]  =  7'b0011101;     //71pi/512
  assign sin[72]  =  7'b1110010;     //72pi/512
  assign cos[72]  =  7'b0011100;     //72pi/512
  assign sin[73]  =  7'b1110010;     //73pi/512
  assign cos[73]  =  7'b0011100;     //73pi/512
  assign sin[74]  =  7'b1110010;     //74pi/512
  assign cos[74]  =  7'b0011100;     //74pi/512
  assign sin[75]  =  7'b1110010;     //75pi/512
  assign cos[75]  =  7'b0011100;     //75pi/512
  assign sin[76]  =  7'b1110010;     //76pi/512
  assign cos[76]  =  7'b0011100;     //76pi/512
  assign sin[77]  =  7'b1110001;     //77pi/512
  assign cos[77]  =  7'b0011100;     //77pi/512
  assign sin[78]  =  7'b1110001;     //78pi/512
  assign cos[78]  =  7'b0011100;     //78pi/512
  assign sin[79]  =  7'b1110001;     //79pi/512
  assign cos[79]  =  7'b0011100;     //79pi/512
  assign sin[80]  =  7'b1110001;     //80pi/512
  assign cos[80]  =  7'b0011100;     //80pi/512
  assign sin[81]  =  7'b1110001;     //81pi/512
  assign cos[81]  =  7'b0011100;     //81pi/512
  assign sin[82]  =  7'b1110001;     //82pi/512
  assign cos[82]  =  7'b0011100;     //82pi/512
  assign sin[83]  =  7'b1110000;     //83pi/512
  assign cos[83]  =  7'b0011011;     //83pi/512
  assign sin[84]  =  7'b1110000;     //84pi/512
  assign cos[84]  =  7'b0011011;     //84pi/512
  assign sin[85]  =  7'b1110000;     //85pi/512
  assign cos[85]  =  7'b0011011;     //85pi/512
  assign sin[86]  =  7'b1110000;     //86pi/512
  assign cos[86]  =  7'b0011011;     //86pi/512
  assign sin[87]  =  7'b1110000;     //87pi/512
  assign cos[87]  =  7'b0011011;     //87pi/512
  assign sin[88]  =  7'b1110000;     //88pi/512
  assign cos[88]  =  7'b0011011;     //88pi/512
  assign sin[89]  =  7'b1101111;     //89pi/512
  assign cos[89]  =  7'b0011011;     //89pi/512
  assign sin[90]  =  7'b1101111;     //90pi/512
  assign cos[90]  =  7'b0011011;     //90pi/512
  assign sin[91]  =  7'b1101111;     //91pi/512
  assign cos[91]  =  7'b0011011;     //91pi/512
  assign sin[92]  =  7'b1101111;     //92pi/512
  assign cos[92]  =  7'b0011011;     //92pi/512
  assign sin[93]  =  7'b1101111;     //93pi/512
  assign cos[93]  =  7'b0011010;     //93pi/512
  assign sin[94]  =  7'b1101111;     //94pi/512
  assign cos[94]  =  7'b0011010;     //94pi/512
  assign sin[95]  =  7'b1101110;     //95pi/512
  assign cos[95]  =  7'b0011010;     //95pi/512
  assign sin[96]  =  7'b1101110;     //96pi/512
  assign cos[96]  =  7'b0011010;     //96pi/512
  assign sin[97]  =  7'b1101110;     //97pi/512
  assign cos[97]  =  7'b0011010;     //97pi/512
  assign sin[98]  =  7'b1101110;     //98pi/512
  assign cos[98]  =  7'b0011010;     //98pi/512
  assign sin[99]  =  7'b1101110;     //99pi/512
  assign cos[99]  =  7'b0011010;     //99pi/512
  assign sin[100]  =  7'b1101110;     //100pi/512
  assign cos[100]  =  7'b0011010;     //100pi/512
  assign sin[101]  =  7'b1101101;     //101pi/512
  assign cos[101]  =  7'b0011010;     //101pi/512
  assign sin[102]  =  7'b1101101;     //102pi/512
  assign cos[102]  =  7'b0011001;     //102pi/512
  assign sin[103]  =  7'b1101101;     //103pi/512
  assign cos[103]  =  7'b0011001;     //103pi/512
  assign sin[104]  =  7'b1101101;     //104pi/512
  assign cos[104]  =  7'b0011001;     //104pi/512
  assign sin[105]  =  7'b1101101;     //105pi/512
  assign cos[105]  =  7'b0011001;     //105pi/512
  assign sin[106]  =  7'b1101101;     //106pi/512
  assign cos[106]  =  7'b0011001;     //106pi/512
  assign sin[107]  =  7'b1101100;     //107pi/512
  assign cos[107]  =  7'b0011001;     //107pi/512
  assign sin[108]  =  7'b1101100;     //108pi/512
  assign cos[108]  =  7'b0011001;     //108pi/512
  assign sin[109]  =  7'b1101100;     //109pi/512
  assign cos[109]  =  7'b0011001;     //109pi/512
  assign sin[110]  =  7'b1101100;     //110pi/512
  assign cos[110]  =  7'b0011000;     //110pi/512
  assign sin[111]  =  7'b1101100;     //111pi/512
  assign cos[111]  =  7'b0011000;     //111pi/512
  assign sin[112]  =  7'b1101100;     //112pi/512
  assign cos[112]  =  7'b0011000;     //112pi/512
  assign sin[113]  =  7'b1101100;     //113pi/512
  assign cos[113]  =  7'b0011000;     //113pi/512
  assign sin[114]  =  7'b1101011;     //114pi/512
  assign cos[114]  =  7'b0011000;     //114pi/512
  assign sin[115]  =  7'b1101011;     //115pi/512
  assign cos[115]  =  7'b0011000;     //115pi/512
  assign sin[116]  =  7'b1101011;     //116pi/512
  assign cos[116]  =  7'b0011000;     //116pi/512
  assign sin[117]  =  7'b1101011;     //117pi/512
  assign cos[117]  =  7'b0011000;     //117pi/512
  assign sin[118]  =  7'b1101011;     //118pi/512
  assign cos[118]  =  7'b0010111;     //118pi/512
  assign sin[119]  =  7'b1101011;     //119pi/512
  assign cos[119]  =  7'b0010111;     //119pi/512
  assign sin[120]  =  7'b1101011;     //120pi/512
  assign cos[120]  =  7'b0010111;     //120pi/512
  assign sin[121]  =  7'b1101010;     //121pi/512
  assign cos[121]  =  7'b0010111;     //121pi/512
  assign sin[122]  =  7'b1101010;     //122pi/512
  assign cos[122]  =  7'b0010111;     //122pi/512
  assign sin[123]  =  7'b1101010;     //123pi/512
  assign cos[123]  =  7'b0010111;     //123pi/512
  assign sin[124]  =  7'b1101010;     //124pi/512
  assign cos[124]  =  7'b0010111;     //124pi/512
  assign sin[125]  =  7'b1101010;     //125pi/512
  assign cos[125]  =  7'b0010111;     //125pi/512
  assign sin[126]  =  7'b1101010;     //126pi/512
  assign cos[126]  =  7'b0010110;     //126pi/512
  assign sin[127]  =  7'b1101010;     //127pi/512
  assign cos[127]  =  7'b0010110;     //127pi/512
  assign sin[128]  =  7'b1101001;     //128pi/512
  assign cos[128]  =  7'b0010110;     //128pi/512
  assign sin[129]  =  7'b1101001;     //129pi/512
  assign cos[129]  =  7'b0010110;     //129pi/512
  assign sin[130]  =  7'b1101001;     //130pi/512
  assign cos[130]  =  7'b0010110;     //130pi/512
  assign sin[131]  =  7'b1101001;     //131pi/512
  assign cos[131]  =  7'b0010110;     //131pi/512
  assign sin[132]  =  7'b1101001;     //132pi/512
  assign cos[132]  =  7'b0010110;     //132pi/512
  assign sin[133]  =  7'b1101001;     //133pi/512
  assign cos[133]  =  7'b0010101;     //133pi/512
  assign sin[134]  =  7'b1101001;     //134pi/512
  assign cos[134]  =  7'b0010101;     //134pi/512
  assign sin[135]  =  7'b1101000;     //135pi/512
  assign cos[135]  =  7'b0010101;     //135pi/512
  assign sin[136]  =  7'b1101000;     //136pi/512
  assign cos[136]  =  7'b0010101;     //136pi/512
  assign sin[137]  =  7'b1101000;     //137pi/512
  assign cos[137]  =  7'b0010101;     //137pi/512
  assign sin[138]  =  7'b1101000;     //138pi/512
  assign cos[138]  =  7'b0010101;     //138pi/512
  assign sin[139]  =  7'b1101000;     //139pi/512
  assign cos[139]  =  7'b0010101;     //139pi/512
  assign sin[140]  =  7'b1101000;     //140pi/512
  assign cos[140]  =  7'b0010100;     //140pi/512
  assign sin[141]  =  7'b1101000;     //141pi/512
  assign cos[141]  =  7'b0010100;     //141pi/512
  assign sin[142]  =  7'b1101000;     //142pi/512
  assign cos[142]  =  7'b0010100;     //142pi/512
  assign sin[143]  =  7'b1100111;     //143pi/512
  assign cos[143]  =  7'b0010100;     //143pi/512
  assign sin[144]  =  7'b1100111;     //144pi/512
  assign cos[144]  =  7'b0010100;     //144pi/512
  assign sin[145]  =  7'b1100111;     //145pi/512
  assign cos[145]  =  7'b0010100;     //145pi/512
  assign sin[146]  =  7'b1100111;     //146pi/512
  assign cos[146]  =  7'b0010011;     //146pi/512
  assign sin[147]  =  7'b1100111;     //147pi/512
  assign cos[147]  =  7'b0010011;     //147pi/512
  assign sin[148]  =  7'b1100111;     //148pi/512
  assign cos[148]  =  7'b0010011;     //148pi/512
  assign sin[149]  =  7'b1100111;     //149pi/512
  assign cos[149]  =  7'b0010011;     //149pi/512
  assign sin[150]  =  7'b1100111;     //150pi/512
  assign cos[150]  =  7'b0010011;     //150pi/512
  assign sin[151]  =  7'b1100110;     //151pi/512
  assign cos[151]  =  7'b0010011;     //151pi/512
  assign sin[152]  =  7'b1100110;     //152pi/512
  assign cos[152]  =  7'b0010011;     //152pi/512
  assign sin[153]  =  7'b1100110;     //153pi/512
  assign cos[153]  =  7'b0010010;     //153pi/512
  assign sin[154]  =  7'b1100110;     //154pi/512
  assign cos[154]  =  7'b0010010;     //154pi/512
  assign sin[155]  =  7'b1100110;     //155pi/512
  assign cos[155]  =  7'b0010010;     //155pi/512
  assign sin[156]  =  7'b1100110;     //156pi/512
  assign cos[156]  =  7'b0010010;     //156pi/512
  assign sin[157]  =  7'b1100110;     //157pi/512
  assign cos[157]  =  7'b0010010;     //157pi/512
  assign sin[158]  =  7'b1100110;     //158pi/512
  assign cos[158]  =  7'b0010010;     //158pi/512
  assign sin[159]  =  7'b1100110;     //159pi/512
  assign cos[159]  =  7'b0010001;     //159pi/512
  assign sin[160]  =  7'b1100101;     //160pi/512
  assign cos[160]  =  7'b0010001;     //160pi/512
  assign sin[161]  =  7'b1100101;     //161pi/512
  assign cos[161]  =  7'b0010001;     //161pi/512
  assign sin[162]  =  7'b1100101;     //162pi/512
  assign cos[162]  =  7'b0010001;     //162pi/512
  assign sin[163]  =  7'b1100101;     //163pi/512
  assign cos[163]  =  7'b0010001;     //163pi/512
  assign sin[164]  =  7'b1100101;     //164pi/512
  assign cos[164]  =  7'b0010001;     //164pi/512
  assign sin[165]  =  7'b1100101;     //165pi/512
  assign cos[165]  =  7'b0010000;     //165pi/512
  assign sin[166]  =  7'b1100101;     //166pi/512
  assign cos[166]  =  7'b0010000;     //166pi/512
  assign sin[167]  =  7'b1100101;     //167pi/512
  assign cos[167]  =  7'b0010000;     //167pi/512
  assign sin[168]  =  7'b1100101;     //168pi/512
  assign cos[168]  =  7'b0010000;     //168pi/512
  assign sin[169]  =  7'b1100100;     //169pi/512
  assign cos[169]  =  7'b0010000;     //169pi/512
  assign sin[170]  =  7'b1100100;     //170pi/512
  assign cos[170]  =  7'b0010000;     //170pi/512
  assign sin[171]  =  7'b1100100;     //171pi/512
  assign cos[171]  =  7'b0001111;     //171pi/512
  assign sin[172]  =  7'b1100100;     //172pi/512
  assign cos[172]  =  7'b0001111;     //172pi/512
  assign sin[173]  =  7'b1100100;     //173pi/512
  assign cos[173]  =  7'b0001111;     //173pi/512
  assign sin[174]  =  7'b1100100;     //174pi/512
  assign cos[174]  =  7'b0001111;     //174pi/512
  assign sin[175]  =  7'b1100100;     //175pi/512
  assign cos[175]  =  7'b0001111;     //175pi/512
  assign sin[176]  =  7'b1100100;     //176pi/512
  assign cos[176]  =  7'b0001111;     //176pi/512
  assign sin[177]  =  7'b1100100;     //177pi/512
  assign cos[177]  =  7'b0001110;     //177pi/512
  assign sin[178]  =  7'b1100100;     //178pi/512
  assign cos[178]  =  7'b0001110;     //178pi/512
  assign sin[179]  =  7'b1100100;     //179pi/512
  assign cos[179]  =  7'b0001110;     //179pi/512
  assign sin[180]  =  7'b1100011;     //180pi/512
  assign cos[180]  =  7'b0001110;     //180pi/512
  assign sin[181]  =  7'b1100011;     //181pi/512
  assign cos[181]  =  7'b0001110;     //181pi/512
  assign sin[182]  =  7'b1100011;     //182pi/512
  assign cos[182]  =  7'b0001110;     //182pi/512
  assign sin[183]  =  7'b1100011;     //183pi/512
  assign cos[183]  =  7'b0001101;     //183pi/512
  assign sin[184]  =  7'b1100011;     //184pi/512
  assign cos[184]  =  7'b0001101;     //184pi/512
  assign sin[185]  =  7'b1100011;     //185pi/512
  assign cos[185]  =  7'b0001101;     //185pi/512
  assign sin[186]  =  7'b1100011;     //186pi/512
  assign cos[186]  =  7'b0001101;     //186pi/512
  assign sin[187]  =  7'b1100011;     //187pi/512
  assign cos[187]  =  7'b0001101;     //187pi/512
  assign sin[188]  =  7'b1100011;     //188pi/512
  assign cos[188]  =  7'b0001100;     //188pi/512
  assign sin[189]  =  7'b1100011;     //189pi/512
  assign cos[189]  =  7'b0001100;     //189pi/512
  assign sin[190]  =  7'b1100011;     //190pi/512
  assign cos[190]  =  7'b0001100;     //190pi/512
  assign sin[191]  =  7'b1100011;     //191pi/512
  assign cos[191]  =  7'b0001100;     //191pi/512
  assign sin[192]  =  7'b1100010;     //192pi/512
  assign cos[192]  =  7'b0001100;     //192pi/512
  assign sin[193]  =  7'b1100010;     //193pi/512
  assign cos[193]  =  7'b0001100;     //193pi/512
  assign sin[194]  =  7'b1100010;     //194pi/512
  assign cos[194]  =  7'b0001011;     //194pi/512
  assign sin[195]  =  7'b1100010;     //195pi/512
  assign cos[195]  =  7'b0001011;     //195pi/512
  assign sin[196]  =  7'b1100010;     //196pi/512
  assign cos[196]  =  7'b0001011;     //196pi/512
  assign sin[197]  =  7'b1100010;     //197pi/512
  assign cos[197]  =  7'b0001011;     //197pi/512
  assign sin[198]  =  7'b1100010;     //198pi/512
  assign cos[198]  =  7'b0001011;     //198pi/512
  assign sin[199]  =  7'b1100010;     //199pi/512
  assign cos[199]  =  7'b0001010;     //199pi/512
  assign sin[200]  =  7'b1100010;     //200pi/512
  assign cos[200]  =  7'b0001010;     //200pi/512
  assign sin[201]  =  7'b1100010;     //201pi/512
  assign cos[201]  =  7'b0001010;     //201pi/512
  assign sin[202]  =  7'b1100010;     //202pi/512
  assign cos[202]  =  7'b0001010;     //202pi/512
  assign sin[203]  =  7'b1100010;     //203pi/512
  assign cos[203]  =  7'b0001010;     //203pi/512
  assign sin[204]  =  7'b1100010;     //204pi/512
  assign cos[204]  =  7'b0001010;     //204pi/512
  assign sin[205]  =  7'b1100010;     //205pi/512
  assign cos[205]  =  7'b0001001;     //205pi/512
  assign sin[206]  =  7'b1100001;     //206pi/512
  assign cos[206]  =  7'b0001001;     //206pi/512
  assign sin[207]  =  7'b1100001;     //207pi/512
  assign cos[207]  =  7'b0001001;     //207pi/512
  assign sin[208]  =  7'b1100001;     //208pi/512
  assign cos[208]  =  7'b0001001;     //208pi/512
  assign sin[209]  =  7'b1100001;     //209pi/512
  assign cos[209]  =  7'b0001001;     //209pi/512
  assign sin[210]  =  7'b1100001;     //210pi/512
  assign cos[210]  =  7'b0001000;     //210pi/512
  assign sin[211]  =  7'b1100001;     //211pi/512
  assign cos[211]  =  7'b0001000;     //211pi/512
  assign sin[212]  =  7'b1100001;     //212pi/512
  assign cos[212]  =  7'b0001000;     //212pi/512
  assign sin[213]  =  7'b1100001;     //213pi/512
  assign cos[213]  =  7'b0001000;     //213pi/512
  assign sin[214]  =  7'b1100001;     //214pi/512
  assign cos[214]  =  7'b0001000;     //214pi/512
  assign sin[215]  =  7'b1100001;     //215pi/512
  assign cos[215]  =  7'b0000111;     //215pi/512
  assign sin[216]  =  7'b1100001;     //216pi/512
  assign cos[216]  =  7'b0000111;     //216pi/512
  assign sin[217]  =  7'b1100001;     //217pi/512
  assign cos[217]  =  7'b0000111;     //217pi/512
  assign sin[218]  =  7'b1100001;     //218pi/512
  assign cos[218]  =  7'b0000111;     //218pi/512
  assign sin[219]  =  7'b1100001;     //219pi/512
  assign cos[219]  =  7'b0000111;     //219pi/512
  assign sin[220]  =  7'b1100001;     //220pi/512
  assign cos[220]  =  7'b0000111;     //220pi/512
  assign sin[221]  =  7'b1100001;     //221pi/512
  assign cos[221]  =  7'b0000110;     //221pi/512
  assign sin[222]  =  7'b1100001;     //222pi/512
  assign cos[222]  =  7'b0000110;     //222pi/512
  assign sin[223]  =  7'b1100001;     //223pi/512
  assign cos[223]  =  7'b0000110;     //223pi/512
  assign sin[224]  =  7'b1100001;     //224pi/512
  assign cos[224]  =  7'b0000110;     //224pi/512
  assign sin[225]  =  7'b1100001;     //225pi/512
  assign cos[225]  =  7'b0000110;     //225pi/512
  assign sin[226]  =  7'b1100001;     //226pi/512
  assign cos[226]  =  7'b0000101;     //226pi/512
  assign sin[227]  =  7'b1100001;     //227pi/512
  assign cos[227]  =  7'b0000101;     //227pi/512
  assign sin[228]  =  7'b1100000;     //228pi/512
  assign cos[228]  =  7'b0000101;     //228pi/512
  assign sin[229]  =  7'b1100000;     //229pi/512
  assign cos[229]  =  7'b0000101;     //229pi/512
  assign sin[230]  =  7'b1100000;     //230pi/512
  assign cos[230]  =  7'b0000101;     //230pi/512
  assign sin[231]  =  7'b1100000;     //231pi/512
  assign cos[231]  =  7'b0000100;     //231pi/512
  assign sin[232]  =  7'b1100000;     //232pi/512
  assign cos[232]  =  7'b0000100;     //232pi/512
  assign sin[233]  =  7'b1100000;     //233pi/512
  assign cos[233]  =  7'b0000100;     //233pi/512
  assign sin[234]  =  7'b1100000;     //234pi/512
  assign cos[234]  =  7'b0000100;     //234pi/512
  assign sin[235]  =  7'b1100000;     //235pi/512
  assign cos[235]  =  7'b0000100;     //235pi/512
  assign sin[236]  =  7'b1100000;     //236pi/512
  assign cos[236]  =  7'b0000011;     //236pi/512
  assign sin[237]  =  7'b1100000;     //237pi/512
  assign cos[237]  =  7'b0000011;     //237pi/512
  assign sin[238]  =  7'b1100000;     //238pi/512
  assign cos[238]  =  7'b0000011;     //238pi/512
  assign sin[239]  =  7'b1100000;     //239pi/512
  assign cos[239]  =  7'b0000011;     //239pi/512
  assign sin[240]  =  7'b1100000;     //240pi/512
  assign cos[240]  =  7'b0000011;     //240pi/512
  assign sin[241]  =  7'b1100000;     //241pi/512
  assign cos[241]  =  7'b0000010;     //241pi/512
  assign sin[242]  =  7'b1100000;     //242pi/512
  assign cos[242]  =  7'b0000010;     //242pi/512
  assign sin[243]  =  7'b1100000;     //243pi/512
  assign cos[243]  =  7'b0000010;     //243pi/512
  assign sin[244]  =  7'b1100000;     //244pi/512
  assign cos[244]  =  7'b0000010;     //244pi/512
  assign sin[245]  =  7'b1100000;     //245pi/512
  assign cos[245]  =  7'b0000010;     //245pi/512
  assign sin[246]  =  7'b1100000;     //246pi/512
  assign cos[246]  =  7'b0000001;     //246pi/512
  assign sin[247]  =  7'b1100000;     //247pi/512
  assign cos[247]  =  7'b0000001;     //247pi/512
  assign sin[248]  =  7'b1100000;     //248pi/512
  assign cos[248]  =  7'b0000001;     //248pi/512
  assign sin[249]  =  7'b1100000;     //249pi/512
  assign cos[249]  =  7'b0000001;     //249pi/512
  assign sin[250]  =  7'b1100000;     //250pi/512
  assign cos[250]  =  7'b0000001;     //250pi/512
  assign sin[251]  =  7'b1100000;     //251pi/512
  assign cos[251]  =  7'b0000000;     //251pi/512
  assign sin[252]  =  7'b1100000;     //252pi/512
  assign cos[252]  =  7'b0000000;     //252pi/512
  assign sin[253]  =  7'b1100000;     //253pi/512
  assign cos[253]  =  7'b0000000;     //253pi/512
  assign sin[254]  =  7'b1100000;     //254pi/512
  assign cos[254]  =  7'b0000000;     //254pi/512
  assign sin[255]  =  7'b1100000;     //255pi/512
  assign cos[255]  =  7'b0000000;     //255pi/512
  assign sin[256]  =  7'b1100000;     //256pi/512
  assign cos[256]  =  7'b0000000;     //256pi/512
  assign sin[257]  =  7'b1100000;     //257pi/512
  assign cos[257]  =  7'b0000000;     //257pi/512
  assign sin[258]  =  7'b1100000;     //258pi/512
  assign cos[258]  =  7'b0000000;     //258pi/512
  assign sin[259]  =  7'b1100000;     //259pi/512
  assign cos[259]  =  7'b1111111;     //259pi/512
  assign sin[260]  =  7'b1100000;     //260pi/512
  assign cos[260]  =  7'b1111111;     //260pi/512
  assign sin[261]  =  7'b1100000;     //261pi/512
  assign cos[261]  =  7'b1111111;     //261pi/512
  assign sin[262]  =  7'b1100000;     //262pi/512
  assign cos[262]  =  7'b1111111;     //262pi/512
  assign sin[263]  =  7'b1100000;     //263pi/512
  assign cos[263]  =  7'b1111111;     //263pi/512
  assign sin[264]  =  7'b1100000;     //264pi/512
  assign cos[264]  =  7'b1111110;     //264pi/512
  assign sin[265]  =  7'b1100000;     //265pi/512
  assign cos[265]  =  7'b1111110;     //265pi/512
  assign sin[266]  =  7'b1100000;     //266pi/512
  assign cos[266]  =  7'b1111110;     //266pi/512
  assign sin[267]  =  7'b1100000;     //267pi/512
  assign cos[267]  =  7'b1111110;     //267pi/512
  assign sin[268]  =  7'b1100000;     //268pi/512
  assign cos[268]  =  7'b1111110;     //268pi/512
  assign sin[269]  =  7'b1100000;     //269pi/512
  assign cos[269]  =  7'b1111101;     //269pi/512
  assign sin[270]  =  7'b1100000;     //270pi/512
  assign cos[270]  =  7'b1111101;     //270pi/512
  assign sin[271]  =  7'b1100000;     //271pi/512
  assign cos[271]  =  7'b1111101;     //271pi/512
  assign sin[272]  =  7'b1100000;     //272pi/512
  assign cos[272]  =  7'b1111101;     //272pi/512
  assign sin[273]  =  7'b1100000;     //273pi/512
  assign cos[273]  =  7'b1111101;     //273pi/512
  assign sin[274]  =  7'b1100000;     //274pi/512
  assign cos[274]  =  7'b1111100;     //274pi/512
  assign sin[275]  =  7'b1100000;     //275pi/512
  assign cos[275]  =  7'b1111100;     //275pi/512
  assign sin[276]  =  7'b1100000;     //276pi/512
  assign cos[276]  =  7'b1111100;     //276pi/512
  assign sin[277]  =  7'b1100000;     //277pi/512
  assign cos[277]  =  7'b1111100;     //277pi/512
  assign sin[278]  =  7'b1100000;     //278pi/512
  assign cos[278]  =  7'b1111100;     //278pi/512
  assign sin[279]  =  7'b1100000;     //279pi/512
  assign cos[279]  =  7'b1111011;     //279pi/512
  assign sin[280]  =  7'b1100000;     //280pi/512
  assign cos[280]  =  7'b1111011;     //280pi/512
  assign sin[281]  =  7'b1100000;     //281pi/512
  assign cos[281]  =  7'b1111011;     //281pi/512
  assign sin[282]  =  7'b1100000;     //282pi/512
  assign cos[282]  =  7'b1111011;     //282pi/512
  assign sin[283]  =  7'b1100000;     //283pi/512
  assign cos[283]  =  7'b1111011;     //283pi/512
  assign sin[284]  =  7'b1100000;     //284pi/512
  assign cos[284]  =  7'b1111011;     //284pi/512
  assign sin[285]  =  7'b1100001;     //285pi/512
  assign cos[285]  =  7'b1111010;     //285pi/512
  assign sin[286]  =  7'b1100001;     //286pi/512
  assign cos[286]  =  7'b1111010;     //286pi/512
  assign sin[287]  =  7'b1100001;     //287pi/512
  assign cos[287]  =  7'b1111010;     //287pi/512
  assign sin[288]  =  7'b1100001;     //288pi/512
  assign cos[288]  =  7'b1111010;     //288pi/512
  assign sin[289]  =  7'b1100001;     //289pi/512
  assign cos[289]  =  7'b1111010;     //289pi/512
  assign sin[290]  =  7'b1100001;     //290pi/512
  assign cos[290]  =  7'b1111001;     //290pi/512
  assign sin[291]  =  7'b1100001;     //291pi/512
  assign cos[291]  =  7'b1111001;     //291pi/512
  assign sin[292]  =  7'b1100001;     //292pi/512
  assign cos[292]  =  7'b1111001;     //292pi/512
  assign sin[293]  =  7'b1100001;     //293pi/512
  assign cos[293]  =  7'b1111001;     //293pi/512
  assign sin[294]  =  7'b1100001;     //294pi/512
  assign cos[294]  =  7'b1111001;     //294pi/512
  assign sin[295]  =  7'b1100001;     //295pi/512
  assign cos[295]  =  7'b1111000;     //295pi/512
  assign sin[296]  =  7'b1100001;     //296pi/512
  assign cos[296]  =  7'b1111000;     //296pi/512
  assign sin[297]  =  7'b1100001;     //297pi/512
  assign cos[297]  =  7'b1111000;     //297pi/512
  assign sin[298]  =  7'b1100001;     //298pi/512
  assign cos[298]  =  7'b1111000;     //298pi/512
  assign sin[299]  =  7'b1100001;     //299pi/512
  assign cos[299]  =  7'b1111000;     //299pi/512
  assign sin[300]  =  7'b1100001;     //300pi/512
  assign cos[300]  =  7'b1110111;     //300pi/512
  assign sin[301]  =  7'b1100001;     //301pi/512
  assign cos[301]  =  7'b1110111;     //301pi/512
  assign sin[302]  =  7'b1100001;     //302pi/512
  assign cos[302]  =  7'b1110111;     //302pi/512
  assign sin[303]  =  7'b1100001;     //303pi/512
  assign cos[303]  =  7'b1110111;     //303pi/512
  assign sin[304]  =  7'b1100001;     //304pi/512
  assign cos[304]  =  7'b1110111;     //304pi/512
  assign sin[305]  =  7'b1100001;     //305pi/512
  assign cos[305]  =  7'b1110111;     //305pi/512
  assign sin[306]  =  7'b1100001;     //306pi/512
  assign cos[306]  =  7'b1110110;     //306pi/512
  assign sin[307]  =  7'b1100010;     //307pi/512
  assign cos[307]  =  7'b1110110;     //307pi/512
  assign sin[308]  =  7'b1100010;     //308pi/512
  assign cos[308]  =  7'b1110110;     //308pi/512
  assign sin[309]  =  7'b1100010;     //309pi/512
  assign cos[309]  =  7'b1110110;     //309pi/512
  assign sin[310]  =  7'b1100010;     //310pi/512
  assign cos[310]  =  7'b1110110;     //310pi/512
  assign sin[311]  =  7'b1100010;     //311pi/512
  assign cos[311]  =  7'b1110101;     //311pi/512
  assign sin[312]  =  7'b1100010;     //312pi/512
  assign cos[312]  =  7'b1110101;     //312pi/512
  assign sin[313]  =  7'b1100010;     //313pi/512
  assign cos[313]  =  7'b1110101;     //313pi/512
  assign sin[314]  =  7'b1100010;     //314pi/512
  assign cos[314]  =  7'b1110101;     //314pi/512
  assign sin[315]  =  7'b1100010;     //315pi/512
  assign cos[315]  =  7'b1110101;     //315pi/512
  assign sin[316]  =  7'b1100010;     //316pi/512
  assign cos[316]  =  7'b1110100;     //316pi/512
  assign sin[317]  =  7'b1100010;     //317pi/512
  assign cos[317]  =  7'b1110100;     //317pi/512
  assign sin[318]  =  7'b1100010;     //318pi/512
  assign cos[318]  =  7'b1110100;     //318pi/512
  assign sin[319]  =  7'b1100010;     //319pi/512
  assign cos[319]  =  7'b1110100;     //319pi/512
  assign sin[320]  =  7'b1100010;     //320pi/512
  assign cos[320]  =  7'b1110100;     //320pi/512
  assign sin[321]  =  7'b1100011;     //321pi/512
  assign cos[321]  =  7'b1110100;     //321pi/512
  assign sin[322]  =  7'b1100011;     //322pi/512
  assign cos[322]  =  7'b1110011;     //322pi/512
  assign sin[323]  =  7'b1100011;     //323pi/512
  assign cos[323]  =  7'b1110011;     //323pi/512
  assign sin[324]  =  7'b1100011;     //324pi/512
  assign cos[324]  =  7'b1110011;     //324pi/512
  assign sin[325]  =  7'b1100011;     //325pi/512
  assign cos[325]  =  7'b1110011;     //325pi/512
  assign sin[326]  =  7'b1100011;     //326pi/512
  assign cos[326]  =  7'b1110011;     //326pi/512
  assign sin[327]  =  7'b1100011;     //327pi/512
  assign cos[327]  =  7'b1110010;     //327pi/512
  assign sin[328]  =  7'b1100011;     //328pi/512
  assign cos[328]  =  7'b1110010;     //328pi/512
  assign sin[329]  =  7'b1100011;     //329pi/512
  assign cos[329]  =  7'b1110010;     //329pi/512
  assign sin[330]  =  7'b1100011;     //330pi/512
  assign cos[330]  =  7'b1110010;     //330pi/512
  assign sin[331]  =  7'b1100011;     //331pi/512
  assign cos[331]  =  7'b1110010;     //331pi/512
  assign sin[332]  =  7'b1100011;     //332pi/512
  assign cos[332]  =  7'b1110010;     //332pi/512
  assign sin[333]  =  7'b1100100;     //333pi/512
  assign cos[333]  =  7'b1110001;     //333pi/512
  assign sin[334]  =  7'b1100100;     //334pi/512
  assign cos[334]  =  7'b1110001;     //334pi/512
  assign sin[335]  =  7'b1100100;     //335pi/512
  assign cos[335]  =  7'b1110001;     //335pi/512
  assign sin[336]  =  7'b1100100;     //336pi/512
  assign cos[336]  =  7'b1110001;     //336pi/512
  assign sin[337]  =  7'b1100100;     //337pi/512
  assign cos[337]  =  7'b1110001;     //337pi/512
  assign sin[338]  =  7'b1100100;     //338pi/512
  assign cos[338]  =  7'b1110001;     //338pi/512
  assign sin[339]  =  7'b1100100;     //339pi/512
  assign cos[339]  =  7'b1110000;     //339pi/512
  assign sin[340]  =  7'b1100100;     //340pi/512
  assign cos[340]  =  7'b1110000;     //340pi/512
  assign sin[341]  =  7'b1100100;     //341pi/512
  assign cos[341]  =  7'b1110000;     //341pi/512
  assign sin[342]  =  7'b1100100;     //342pi/512
  assign cos[342]  =  7'b1110000;     //342pi/512
  assign sin[343]  =  7'b1100100;     //343pi/512
  assign cos[343]  =  7'b1110000;     //343pi/512
  assign sin[344]  =  7'b1100101;     //344pi/512
  assign cos[344]  =  7'b1110000;     //344pi/512
  assign sin[345]  =  7'b1100101;     //345pi/512
  assign cos[345]  =  7'b1101111;     //345pi/512
  assign sin[346]  =  7'b1100101;     //346pi/512
  assign cos[346]  =  7'b1101111;     //346pi/512
  assign sin[347]  =  7'b1100101;     //347pi/512
  assign cos[347]  =  7'b1101111;     //347pi/512
  assign sin[348]  =  7'b1100101;     //348pi/512
  assign cos[348]  =  7'b1101111;     //348pi/512
  assign sin[349]  =  7'b1100101;     //349pi/512
  assign cos[349]  =  7'b1101111;     //349pi/512
  assign sin[350]  =  7'b1100101;     //350pi/512
  assign cos[350]  =  7'b1101111;     //350pi/512
  assign sin[351]  =  7'b1100101;     //351pi/512
  assign cos[351]  =  7'b1101110;     //351pi/512
  assign sin[352]  =  7'b1100101;     //352pi/512
  assign cos[352]  =  7'b1101110;     //352pi/512
  assign sin[353]  =  7'b1100110;     //353pi/512
  assign cos[353]  =  7'b1101110;     //353pi/512
  assign sin[354]  =  7'b1100110;     //354pi/512
  assign cos[354]  =  7'b1101110;     //354pi/512
  assign sin[355]  =  7'b1100110;     //355pi/512
  assign cos[355]  =  7'b1101110;     //355pi/512
  assign sin[356]  =  7'b1100110;     //356pi/512
  assign cos[356]  =  7'b1101110;     //356pi/512
  assign sin[357]  =  7'b1100110;     //357pi/512
  assign cos[357]  =  7'b1101101;     //357pi/512
  assign sin[358]  =  7'b1100110;     //358pi/512
  assign cos[358]  =  7'b1101101;     //358pi/512
  assign sin[359]  =  7'b1100110;     //359pi/512
  assign cos[359]  =  7'b1101101;     //359pi/512
  assign sin[360]  =  7'b1100110;     //360pi/512
  assign cos[360]  =  7'b1101101;     //360pi/512
  assign sin[361]  =  7'b1100110;     //361pi/512
  assign cos[361]  =  7'b1101101;     //361pi/512
  assign sin[362]  =  7'b1100111;     //362pi/512
  assign cos[362]  =  7'b1101101;     //362pi/512
  assign sin[363]  =  7'b1100111;     //363pi/512
  assign cos[363]  =  7'b1101100;     //363pi/512
  assign sin[364]  =  7'b1100111;     //364pi/512
  assign cos[364]  =  7'b1101100;     //364pi/512
  assign sin[365]  =  7'b1100111;     //365pi/512
  assign cos[365]  =  7'b1101100;     //365pi/512
  assign sin[366]  =  7'b1100111;     //366pi/512
  assign cos[366]  =  7'b1101100;     //366pi/512
  assign sin[367]  =  7'b1100111;     //367pi/512
  assign cos[367]  =  7'b1101100;     //367pi/512
  assign sin[368]  =  7'b1100111;     //368pi/512
  assign cos[368]  =  7'b1101100;     //368pi/512
  assign sin[369]  =  7'b1100111;     //369pi/512
  assign cos[369]  =  7'b1101100;     //369pi/512
  assign sin[370]  =  7'b1101000;     //370pi/512
  assign cos[370]  =  7'b1101011;     //370pi/512
  assign sin[371]  =  7'b1101000;     //371pi/512
  assign cos[371]  =  7'b1101011;     //371pi/512
  assign sin[372]  =  7'b1101000;     //372pi/512
  assign cos[372]  =  7'b1101011;     //372pi/512
  assign sin[373]  =  7'b1101000;     //373pi/512
  assign cos[373]  =  7'b1101011;     //373pi/512
  assign sin[374]  =  7'b1101000;     //374pi/512
  assign cos[374]  =  7'b1101011;     //374pi/512
  assign sin[375]  =  7'b1101000;     //375pi/512
  assign cos[375]  =  7'b1101011;     //375pi/512
  assign sin[376]  =  7'b1101000;     //376pi/512
  assign cos[376]  =  7'b1101011;     //376pi/512
  assign sin[377]  =  7'b1101000;     //377pi/512
  assign cos[377]  =  7'b1101010;     //377pi/512
  assign sin[378]  =  7'b1101001;     //378pi/512
  assign cos[378]  =  7'b1101010;     //378pi/512
  assign sin[379]  =  7'b1101001;     //379pi/512
  assign cos[379]  =  7'b1101010;     //379pi/512
  assign sin[380]  =  7'b1101001;     //380pi/512
  assign cos[380]  =  7'b1101010;     //380pi/512
  assign sin[381]  =  7'b1101001;     //381pi/512
  assign cos[381]  =  7'b1101010;     //381pi/512
  assign sin[382]  =  7'b1101001;     //382pi/512
  assign cos[382]  =  7'b1101010;     //382pi/512
  assign sin[383]  =  7'b1101001;     //383pi/512
  assign cos[383]  =  7'b1101010;     //383pi/512
  assign sin[384]  =  7'b1101001;     //384pi/512
  assign cos[384]  =  7'b1101001;     //384pi/512
  assign sin[385]  =  7'b1101010;     //385pi/512
  assign cos[385]  =  7'b1101001;     //385pi/512
  assign sin[386]  =  7'b1101010;     //386pi/512
  assign cos[386]  =  7'b1101001;     //386pi/512
  assign sin[387]  =  7'b1101010;     //387pi/512
  assign cos[387]  =  7'b1101001;     //387pi/512
  assign sin[388]  =  7'b1101010;     //388pi/512
  assign cos[388]  =  7'b1101001;     //388pi/512
  assign sin[389]  =  7'b1101010;     //389pi/512
  assign cos[389]  =  7'b1101001;     //389pi/512
  assign sin[390]  =  7'b1101010;     //390pi/512
  assign cos[390]  =  7'b1101001;     //390pi/512
  assign sin[391]  =  7'b1101010;     //391pi/512
  assign cos[391]  =  7'b1101000;     //391pi/512
  assign sin[392]  =  7'b1101011;     //392pi/512
  assign cos[392]  =  7'b1101000;     //392pi/512
  assign sin[393]  =  7'b1101011;     //393pi/512
  assign cos[393]  =  7'b1101000;     //393pi/512
  assign sin[394]  =  7'b1101011;     //394pi/512
  assign cos[394]  =  7'b1101000;     //394pi/512
  assign sin[395]  =  7'b1101011;     //395pi/512
  assign cos[395]  =  7'b1101000;     //395pi/512
  assign sin[396]  =  7'b1101011;     //396pi/512
  assign cos[396]  =  7'b1101000;     //396pi/512
  assign sin[397]  =  7'b1101011;     //397pi/512
  assign cos[397]  =  7'b1101000;     //397pi/512
  assign sin[398]  =  7'b1101011;     //398pi/512
  assign cos[398]  =  7'b1101000;     //398pi/512
  assign sin[399]  =  7'b1101100;     //399pi/512
  assign cos[399]  =  7'b1100111;     //399pi/512
  assign sin[400]  =  7'b1101100;     //400pi/512
  assign cos[400]  =  7'b1100111;     //400pi/512
  assign sin[401]  =  7'b1101100;     //401pi/512
  assign cos[401]  =  7'b1100111;     //401pi/512
  assign sin[402]  =  7'b1101100;     //402pi/512
  assign cos[402]  =  7'b1100111;     //402pi/512
  assign sin[403]  =  7'b1101100;     //403pi/512
  assign cos[403]  =  7'b1100111;     //403pi/512
  assign sin[404]  =  7'b1101100;     //404pi/512
  assign cos[404]  =  7'b1100111;     //404pi/512
  assign sin[405]  =  7'b1101100;     //405pi/512
  assign cos[405]  =  7'b1100111;     //405pi/512
  assign sin[406]  =  7'b1101101;     //406pi/512
  assign cos[406]  =  7'b1100111;     //406pi/512
  assign sin[407]  =  7'b1101101;     //407pi/512
  assign cos[407]  =  7'b1100110;     //407pi/512
  assign sin[408]  =  7'b1101101;     //408pi/512
  assign cos[408]  =  7'b1100110;     //408pi/512
  assign sin[409]  =  7'b1101101;     //409pi/512
  assign cos[409]  =  7'b1100110;     //409pi/512
  assign sin[410]  =  7'b1101101;     //410pi/512
  assign cos[410]  =  7'b1100110;     //410pi/512
  assign sin[411]  =  7'b1101101;     //411pi/512
  assign cos[411]  =  7'b1100110;     //411pi/512
  assign sin[412]  =  7'b1101110;     //412pi/512
  assign cos[412]  =  7'b1100110;     //412pi/512
  assign sin[413]  =  7'b1101110;     //413pi/512
  assign cos[413]  =  7'b1100110;     //413pi/512
  assign sin[414]  =  7'b1101110;     //414pi/512
  assign cos[414]  =  7'b1100110;     //414pi/512
  assign sin[415]  =  7'b1101110;     //415pi/512
  assign cos[415]  =  7'b1100110;     //415pi/512
  assign sin[416]  =  7'b1101110;     //416pi/512
  assign cos[416]  =  7'b1100101;     //416pi/512
  assign sin[417]  =  7'b1101110;     //417pi/512
  assign cos[417]  =  7'b1100101;     //417pi/512
  assign sin[418]  =  7'b1101111;     //418pi/512
  assign cos[418]  =  7'b1100101;     //418pi/512
  assign sin[419]  =  7'b1101111;     //419pi/512
  assign cos[419]  =  7'b1100101;     //419pi/512
  assign sin[420]  =  7'b1101111;     //420pi/512
  assign cos[420]  =  7'b1100101;     //420pi/512
  assign sin[421]  =  7'b1101111;     //421pi/512
  assign cos[421]  =  7'b1100101;     //421pi/512
  assign sin[422]  =  7'b1101111;     //422pi/512
  assign cos[422]  =  7'b1100101;     //422pi/512
  assign sin[423]  =  7'b1101111;     //423pi/512
  assign cos[423]  =  7'b1100101;     //423pi/512
  assign sin[424]  =  7'b1110000;     //424pi/512
  assign cos[424]  =  7'b1100101;     //424pi/512
  assign sin[425]  =  7'b1110000;     //425pi/512
  assign cos[425]  =  7'b1100100;     //425pi/512
  assign sin[426]  =  7'b1110000;     //426pi/512
  assign cos[426]  =  7'b1100100;     //426pi/512
  assign sin[427]  =  7'b1110000;     //427pi/512
  assign cos[427]  =  7'b1100100;     //427pi/512
  assign sin[428]  =  7'b1110000;     //428pi/512
  assign cos[428]  =  7'b1100100;     //428pi/512
  assign sin[429]  =  7'b1110000;     //429pi/512
  assign cos[429]  =  7'b1100100;     //429pi/512
  assign sin[430]  =  7'b1110001;     //430pi/512
  assign cos[430]  =  7'b1100100;     //430pi/512
  assign sin[431]  =  7'b1110001;     //431pi/512
  assign cos[431]  =  7'b1100100;     //431pi/512
  assign sin[432]  =  7'b1110001;     //432pi/512
  assign cos[432]  =  7'b1100100;     //432pi/512
  assign sin[433]  =  7'b1110001;     //433pi/512
  assign cos[433]  =  7'b1100100;     //433pi/512
  assign sin[434]  =  7'b1110001;     //434pi/512
  assign cos[434]  =  7'b1100100;     //434pi/512
  assign sin[435]  =  7'b1110001;     //435pi/512
  assign cos[435]  =  7'b1100100;     //435pi/512
  assign sin[436]  =  7'b1110010;     //436pi/512
  assign cos[436]  =  7'b1100011;     //436pi/512
  assign sin[437]  =  7'b1110010;     //437pi/512
  assign cos[437]  =  7'b1100011;     //437pi/512
  assign sin[438]  =  7'b1110010;     //438pi/512
  assign cos[438]  =  7'b1100011;     //438pi/512
  assign sin[439]  =  7'b1110010;     //439pi/512
  assign cos[439]  =  7'b1100011;     //439pi/512
  assign sin[440]  =  7'b1110010;     //440pi/512
  assign cos[440]  =  7'b1100011;     //440pi/512
  assign sin[441]  =  7'b1110010;     //441pi/512
  assign cos[441]  =  7'b1100011;     //441pi/512
  assign sin[442]  =  7'b1110011;     //442pi/512
  assign cos[442]  =  7'b1100011;     //442pi/512
  assign sin[443]  =  7'b1110011;     //443pi/512
  assign cos[443]  =  7'b1100011;     //443pi/512
  assign sin[444]  =  7'b1110011;     //444pi/512
  assign cos[444]  =  7'b1100011;     //444pi/512
  assign sin[445]  =  7'b1110011;     //445pi/512
  assign cos[445]  =  7'b1100011;     //445pi/512
  assign sin[446]  =  7'b1110011;     //446pi/512
  assign cos[446]  =  7'b1100011;     //446pi/512
  assign sin[447]  =  7'b1110100;     //447pi/512
  assign cos[447]  =  7'b1100011;     //447pi/512
  assign sin[448]  =  7'b1110100;     //448pi/512
  assign cos[448]  =  7'b1100010;     //448pi/512
  assign sin[449]  =  7'b1110100;     //449pi/512
  assign cos[449]  =  7'b1100010;     //449pi/512
  assign sin[450]  =  7'b1110100;     //450pi/512
  assign cos[450]  =  7'b1100010;     //450pi/512
  assign sin[451]  =  7'b1110100;     //451pi/512
  assign cos[451]  =  7'b1100010;     //451pi/512
  assign sin[452]  =  7'b1110100;     //452pi/512
  assign cos[452]  =  7'b1100010;     //452pi/512
  assign sin[453]  =  7'b1110101;     //453pi/512
  assign cos[453]  =  7'b1100010;     //453pi/512
  assign sin[454]  =  7'b1110101;     //454pi/512
  assign cos[454]  =  7'b1100010;     //454pi/512
  assign sin[455]  =  7'b1110101;     //455pi/512
  assign cos[455]  =  7'b1100010;     //455pi/512
  assign sin[456]  =  7'b1110101;     //456pi/512
  assign cos[456]  =  7'b1100010;     //456pi/512
  assign sin[457]  =  7'b1110101;     //457pi/512
  assign cos[457]  =  7'b1100010;     //457pi/512
  assign sin[458]  =  7'b1110110;     //458pi/512
  assign cos[458]  =  7'b1100010;     //458pi/512
  assign sin[459]  =  7'b1110110;     //459pi/512
  assign cos[459]  =  7'b1100010;     //459pi/512
  assign sin[460]  =  7'b1110110;     //460pi/512
  assign cos[460]  =  7'b1100010;     //460pi/512
  assign sin[461]  =  7'b1110110;     //461pi/512
  assign cos[461]  =  7'b1100010;     //461pi/512
  assign sin[462]  =  7'b1110110;     //462pi/512
  assign cos[462]  =  7'b1100001;     //462pi/512
  assign sin[463]  =  7'b1110111;     //463pi/512
  assign cos[463]  =  7'b1100001;     //463pi/512
  assign sin[464]  =  7'b1110111;     //464pi/512
  assign cos[464]  =  7'b1100001;     //464pi/512
  assign sin[465]  =  7'b1110111;     //465pi/512
  assign cos[465]  =  7'b1100001;     //465pi/512
  assign sin[466]  =  7'b1110111;     //466pi/512
  assign cos[466]  =  7'b1100001;     //466pi/512
  assign sin[467]  =  7'b1110111;     //467pi/512
  assign cos[467]  =  7'b1100001;     //467pi/512
  assign sin[468]  =  7'b1110111;     //468pi/512
  assign cos[468]  =  7'b1100001;     //468pi/512
  assign sin[469]  =  7'b1111000;     //469pi/512
  assign cos[469]  =  7'b1100001;     //469pi/512
  assign sin[470]  =  7'b1111000;     //470pi/512
  assign cos[470]  =  7'b1100001;     //470pi/512
  assign sin[471]  =  7'b1111000;     //471pi/512
  assign cos[471]  =  7'b1100001;     //471pi/512
  assign sin[472]  =  7'b1111000;     //472pi/512
  assign cos[472]  =  7'b1100001;     //472pi/512
  assign sin[473]  =  7'b1111000;     //473pi/512
  assign cos[473]  =  7'b1100001;     //473pi/512
  assign sin[474]  =  7'b1111001;     //474pi/512
  assign cos[474]  =  7'b1100001;     //474pi/512
  assign sin[475]  =  7'b1111001;     //475pi/512
  assign cos[475]  =  7'b1100001;     //475pi/512
  assign sin[476]  =  7'b1111001;     //476pi/512
  assign cos[476]  =  7'b1100001;     //476pi/512
  assign sin[477]  =  7'b1111001;     //477pi/512
  assign cos[477]  =  7'b1100001;     //477pi/512
  assign sin[478]  =  7'b1111001;     //478pi/512
  assign cos[478]  =  7'b1100001;     //478pi/512
  assign sin[479]  =  7'b1111010;     //479pi/512
  assign cos[479]  =  7'b1100001;     //479pi/512
  assign sin[480]  =  7'b1111010;     //480pi/512
  assign cos[480]  =  7'b1100001;     //480pi/512
  assign sin[481]  =  7'b1111010;     //481pi/512
  assign cos[481]  =  7'b1100001;     //481pi/512
  assign sin[482]  =  7'b1111010;     //482pi/512
  assign cos[482]  =  7'b1100001;     //482pi/512
  assign sin[483]  =  7'b1111010;     //483pi/512
  assign cos[483]  =  7'b1100001;     //483pi/512
  assign sin[484]  =  7'b1111011;     //484pi/512
  assign cos[484]  =  7'b1100000;     //484pi/512
  assign sin[485]  =  7'b1111011;     //485pi/512
  assign cos[485]  =  7'b1100000;     //485pi/512
  assign sin[486]  =  7'b1111011;     //486pi/512
  assign cos[486]  =  7'b1100000;     //486pi/512
  assign sin[487]  =  7'b1111011;     //487pi/512
  assign cos[487]  =  7'b1100000;     //487pi/512
  assign sin[488]  =  7'b1111011;     //488pi/512
  assign cos[488]  =  7'b1100000;     //488pi/512
  assign sin[489]  =  7'b1111011;     //489pi/512
  assign cos[489]  =  7'b1100000;     //489pi/512
  assign sin[490]  =  7'b1111100;     //490pi/512
  assign cos[490]  =  7'b1100000;     //490pi/512
  assign sin[491]  =  7'b1111100;     //491pi/512
  assign cos[491]  =  7'b1100000;     //491pi/512
  assign sin[492]  =  7'b1111100;     //492pi/512
  assign cos[492]  =  7'b1100000;     //492pi/512
  assign sin[493]  =  7'b1111100;     //493pi/512
  assign cos[493]  =  7'b1100000;     //493pi/512
  assign sin[494]  =  7'b1111100;     //494pi/512
  assign cos[494]  =  7'b1100000;     //494pi/512
  assign sin[495]  =  7'b1111101;     //495pi/512
  assign cos[495]  =  7'b1100000;     //495pi/512
  assign sin[496]  =  7'b1111101;     //496pi/512
  assign cos[496]  =  7'b1100000;     //496pi/512
  assign sin[497]  =  7'b1111101;     //497pi/512
  assign cos[497]  =  7'b1100000;     //497pi/512
  assign sin[498]  =  7'b1111101;     //498pi/512
  assign cos[498]  =  7'b1100000;     //498pi/512
  assign sin[499]  =  7'b1111101;     //499pi/512
  assign cos[499]  =  7'b1100000;     //499pi/512
  assign sin[500]  =  7'b1111110;     //500pi/512
  assign cos[500]  =  7'b1100000;     //500pi/512
  assign sin[501]  =  7'b1111110;     //501pi/512
  assign cos[501]  =  7'b1100000;     //501pi/512
  assign sin[502]  =  7'b1111110;     //502pi/512
  assign cos[502]  =  7'b1100000;     //502pi/512
  assign sin[503]  =  7'b1111110;     //503pi/512
  assign cos[503]  =  7'b1100000;     //503pi/512
  assign sin[504]  =  7'b1111110;     //504pi/512
  assign cos[504]  =  7'b1100000;     //504pi/512
  assign sin[505]  =  7'b1111111;     //505pi/512
  assign cos[505]  =  7'b1100000;     //505pi/512
  assign sin[506]  =  7'b1111111;     //506pi/512
  assign cos[506]  =  7'b1100000;     //506pi/512
  assign sin[507]  =  7'b1111111;     //507pi/512
  assign cos[507]  =  7'b1100000;     //507pi/512
  assign sin[508]  =  7'b1111111;     //508pi/512
  assign cos[508]  =  7'b1100000;     //508pi/512
  assign sin[509]  =  7'b1111111;     //509pi/512
  assign cos[509]  =  7'b1100000;     //509pi/512
  assign sin[510]  =  7'b0000000;     //510pi/512
  assign cos[510]  =  7'b1100000;     //510pi/512
  assign sin[511]  =  7'b0000000;     //511pi/512
  assign cos[511]  =  7'b1100000;     //511pi/512

  ////////////////////////////////////////////////////////
    assign sin2[0]  =  7'b0000000;     //0pi/512
  assign cos2[0]  =  7'b0100000;     //0pi/512
  assign sin2[1]  =  7'b0000000;     //1pi/512
  assign cos2[1]  =  7'b0011111;     //1pi/512
  assign sin2[2]  =  7'b0000000;     //2pi/512
  assign cos2[2]  =  7'b0011111;     //2pi/512
  assign sin2[3]  =  7'b0000000;     //3pi/512
  assign cos2[3]  =  7'b0011111;     //3pi/512
  assign sin2[4]  =  7'b1111111;     //4pi/512
  assign cos2[4]  =  7'b0011111;     //4pi/512
  assign sin2[5]  =  7'b1111111;     //5pi/512
  assign cos2[5]  =  7'b0011111;     //5pi/512
  assign sin2[6]  =  7'b1111111;     //6pi/512
  assign cos2[6]  =  7'b0011111;     //6pi/512
  assign sin2[7]  =  7'b1111111;     //7pi/512
  assign cos2[7]  =  7'b0011111;     //7pi/512
  assign sin2[8]  =  7'b1111111;     //8pi/512
  assign cos2[8]  =  7'b0011111;     //8pi/512
  assign sin2[9]  =  7'b1111111;     //9pi/512
  assign cos2[9]  =  7'b0011111;     //9pi/512
  assign sin2[10]  =  7'b1111110;     //10pi/512
  assign cos2[10]  =  7'b0011111;     //10pi/512
  assign sin2[11]  =  7'b1111110;     //11pi/512
  assign cos2[11]  =  7'b0011111;     //11pi/512
  assign sin2[12]  =  7'b1111110;     //12pi/512
  assign cos2[12]  =  7'b0011111;     //12pi/512
  assign sin2[13]  =  7'b1111110;     //13pi/512
  assign cos2[13]  =  7'b0011111;     //13pi/512
  assign sin2[14]  =  7'b1111110;     //14pi/512
  assign cos2[14]  =  7'b0011111;     //14pi/512
  assign sin2[15]  =  7'b1111110;     //15pi/512
  assign cos2[15]  =  7'b0011111;     //15pi/512
  assign sin2[16]  =  7'b1111101;     //16pi/512
  assign cos2[16]  =  7'b0011111;     //16pi/512
  assign sin2[17]  =  7'b1111101;     //17pi/512
  assign cos2[17]  =  7'b0011111;     //17pi/512
  assign sin2[18]  =  7'b1111101;     //18pi/512
  assign cos2[18]  =  7'b0011111;     //18pi/512
  assign sin2[19]  =  7'b1111101;     //19pi/512
  assign cos2[19]  =  7'b0011111;     //19pi/512
  assign sin2[20]  =  7'b1111101;     //20pi/512
  assign cos2[20]  =  7'b0011111;     //20pi/512
  assign sin2[21]  =  7'b1111101;     //21pi/512
  assign cos2[21]  =  7'b0011111;     //21pi/512
  assign sin2[22]  =  7'b1111101;     //22pi/512
  assign cos2[22]  =  7'b0011111;     //22pi/512
  assign sin2[23]  =  7'b1111100;     //23pi/512
  assign cos2[23]  =  7'b0011111;     //23pi/512
  assign sin2[24]  =  7'b1111100;     //24pi/512
  assign cos2[24]  =  7'b0011111;     //24pi/512
  assign sin2[25]  =  7'b1111100;     //25pi/512
  assign cos2[25]  =  7'b0011111;     //25pi/512
  assign sin2[26]  =  7'b1111100;     //26pi/512
  assign cos2[26]  =  7'b0011111;     //26pi/512
  assign sin2[27]  =  7'b1111100;     //27pi/512
  assign cos2[27]  =  7'b0011111;     //27pi/512
  assign sin2[28]  =  7'b1111100;     //28pi/512
  assign cos2[28]  =  7'b0011111;     //28pi/512
  assign sin2[29]  =  7'b1111011;     //29pi/512
  assign cos2[29]  =  7'b0011111;     //29pi/512
  assign sin2[30]  =  7'b1111011;     //30pi/512
  assign cos2[30]  =  7'b0011111;     //30pi/512
  assign sin2[31]  =  7'b1111011;     //31pi/512
  assign cos2[31]  =  7'b0011111;     //31pi/512
  assign sin2[32]  =  7'b1111011;     //32pi/512
  assign cos2[32]  =  7'b0011111;     //32pi/512
  assign sin2[33]  =  7'b1111011;     //33pi/512
  assign cos2[33]  =  7'b0011111;     //33pi/512
  assign sin2[34]  =  7'b1111011;     //34pi/512
  assign cos2[34]  =  7'b0011111;     //34pi/512
  assign sin2[35]  =  7'b1111011;     //35pi/512
  assign cos2[35]  =  7'b0011111;     //35pi/512
  assign sin2[36]  =  7'b1111010;     //36pi/512
  assign cos2[36]  =  7'b0011111;     //36pi/512
  assign sin2[37]  =  7'b1111010;     //37pi/512
  assign cos2[37]  =  7'b0011111;     //37pi/512
  assign sin2[38]  =  7'b1111010;     //38pi/512
  assign cos2[38]  =  7'b0011111;     //38pi/512
  assign sin2[39]  =  7'b1111010;     //39pi/512
  assign cos2[39]  =  7'b0011111;     //39pi/512
  assign sin2[40]  =  7'b1111010;     //40pi/512
  assign cos2[40]  =  7'b0011111;     //40pi/512
  assign sin2[41]  =  7'b1111010;     //41pi/512
  assign cos2[41]  =  7'b0011111;     //41pi/512
  assign sin2[42]  =  7'b1111001;     //42pi/512
  assign cos2[42]  =  7'b0011111;     //42pi/512
  assign sin2[43]  =  7'b1111001;     //43pi/512
  assign cos2[43]  =  7'b0011111;     //43pi/512
  assign sin2[44]  =  7'b1111001;     //44pi/512
  assign cos2[44]  =  7'b0011111;     //44pi/512
  assign sin2[45]  =  7'b1111001;     //45pi/512
  assign cos2[45]  =  7'b0011111;     //45pi/512
  assign sin2[46]  =  7'b1111001;     //46pi/512
  assign cos2[46]  =  7'b0011111;     //46pi/512
  assign sin2[47]  =  7'b1111001;     //47pi/512
  assign cos2[47]  =  7'b0011111;     //47pi/512
  assign sin2[48]  =  7'b1111001;     //48pi/512
  assign cos2[48]  =  7'b0011111;     //48pi/512
  assign sin2[49]  =  7'b1111000;     //49pi/512
  assign cos2[49]  =  7'b0011111;     //49pi/512
  assign sin2[50]  =  7'b1111000;     //50pi/512
  assign cos2[50]  =  7'b0011111;     //50pi/512
  assign sin2[51]  =  7'b1111000;     //51pi/512
  assign cos2[51]  =  7'b0011111;     //51pi/512
  assign sin2[52]  =  7'b1111000;     //52pi/512
  assign cos2[52]  =  7'b0011110;     //52pi/512
  assign sin2[53]  =  7'b1111000;     //53pi/512
  assign cos2[53]  =  7'b0011110;     //53pi/512
  assign sin2[54]  =  7'b1111000;     //54pi/512
  assign cos2[54]  =  7'b0011110;     //54pi/512
  assign sin2[55]  =  7'b1110111;     //55pi/512
  assign cos2[55]  =  7'b0011110;     //55pi/512
  assign sin2[56]  =  7'b1110111;     //56pi/512
  assign cos2[56]  =  7'b0011110;     //56pi/512
  assign sin2[57]  =  7'b1110111;     //57pi/512
  assign cos2[57]  =  7'b0011110;     //57pi/512
  assign sin2[58]  =  7'b1110111;     //58pi/512
  assign cos2[58]  =  7'b0011110;     //58pi/512
  assign sin2[59]  =  7'b1110111;     //59pi/512
  assign cos2[59]  =  7'b0011110;     //59pi/512
  assign sin2[60]  =  7'b1110111;     //60pi/512
  assign cos2[60]  =  7'b0011110;     //60pi/512
  assign sin2[61]  =  7'b1110111;     //61pi/512
  assign cos2[61]  =  7'b0011110;     //61pi/512
  assign sin2[62]  =  7'b1110110;     //62pi/512
  assign cos2[62]  =  7'b0011110;     //62pi/512
  assign sin2[63]  =  7'b1110110;     //63pi/512
  assign cos2[63]  =  7'b0011110;     //63pi/512
  assign sin2[64]  =  7'b1110110;     //64pi/512
  assign cos2[64]  =  7'b0011110;     //64pi/512
  assign sin2[65]  =  7'b1110110;     //65pi/512
  assign cos2[65]  =  7'b0011110;     //65pi/512
  assign sin2[66]  =  7'b1110110;     //66pi/512
  assign cos2[66]  =  7'b0011110;     //66pi/512
  assign sin2[67]  =  7'b1110110;     //67pi/512
  assign cos2[67]  =  7'b0011110;     //67pi/512
  assign sin2[68]  =  7'b1110110;     //68pi/512
  assign cos2[68]  =  7'b0011110;     //68pi/512
  assign sin2[69]  =  7'b1110101;     //69pi/512
  assign cos2[69]  =  7'b0011110;     //69pi/512
  assign sin2[70]  =  7'b1110101;     //70pi/512
  assign cos2[70]  =  7'b0011110;     //70pi/512
  assign sin2[71]  =  7'b1110101;     //71pi/512
  assign cos2[71]  =  7'b0011110;     //71pi/512
  assign sin2[72]  =  7'b1110101;     //72pi/512
  assign cos2[72]  =  7'b0011110;     //72pi/512
  assign sin2[73]  =  7'b1110101;     //73pi/512
  assign cos2[73]  =  7'b0011101;     //73pi/512
  assign sin2[74]  =  7'b1110101;     //74pi/512
  assign cos2[74]  =  7'b0011101;     //74pi/512
  assign sin2[75]  =  7'b1110100;     //75pi/512
  assign cos2[75]  =  7'b0011101;     //75pi/512
  assign sin2[76]  =  7'b1110100;     //76pi/512
  assign cos2[76]  =  7'b0011101;     //76pi/512
  assign sin2[77]  =  7'b1110100;     //77pi/512
  assign cos2[77]  =  7'b0011101;     //77pi/512
  assign sin2[78]  =  7'b1110100;     //78pi/512
  assign cos2[78]  =  7'b0011101;     //78pi/512
  assign sin2[79]  =  7'b1110100;     //79pi/512
  assign cos2[79]  =  7'b0011101;     //79pi/512
  assign sin2[80]  =  7'b1110100;     //80pi/512
  assign cos2[80]  =  7'b0011101;     //80pi/512
  assign sin2[81]  =  7'b1110100;     //81pi/512
  assign cos2[81]  =  7'b0011101;     //81pi/512
  assign sin2[82]  =  7'b1110011;     //82pi/512
  assign cos2[82]  =  7'b0011101;     //82pi/512
  assign sin2[83]  =  7'b1110011;     //83pi/512
  assign cos2[83]  =  7'b0011101;     //83pi/512
  assign sin2[84]  =  7'b1110011;     //84pi/512
  assign cos2[84]  =  7'b0011101;     //84pi/512
  assign sin2[85]  =  7'b1110011;     //85pi/512
  assign cos2[85]  =  7'b0011101;     //85pi/512
  assign sin2[86]  =  7'b1110011;     //86pi/512
  assign cos2[86]  =  7'b0011101;     //86pi/512
  assign sin2[87]  =  7'b1110011;     //87pi/512
  assign cos2[87]  =  7'b0011101;     //87pi/512
  assign sin2[88]  =  7'b1110011;     //88pi/512
  assign cos2[88]  =  7'b0011101;     //88pi/512
  assign sin2[89]  =  7'b1110010;     //89pi/512
  assign cos2[89]  =  7'b0011100;     //89pi/512
  assign sin2[90]  =  7'b1110010;     //90pi/512
  assign cos2[90]  =  7'b0011100;     //90pi/512
  assign sin2[91]  =  7'b1110010;     //91pi/512
  assign cos2[91]  =  7'b0011100;     //91pi/512
  assign sin2[92]  =  7'b1110010;     //92pi/512
  assign cos2[92]  =  7'b0011100;     //92pi/512
  assign sin2[93]  =  7'b1110010;     //93pi/512
  assign cos2[93]  =  7'b0011100;     //93pi/512
  assign sin2[94]  =  7'b1110010;     //94pi/512
  assign cos2[94]  =  7'b0011100;     //94pi/512
  assign sin2[95]  =  7'b1110010;     //95pi/512
  assign cos2[95]  =  7'b0011100;     //95pi/512
  assign sin2[96]  =  7'b1110001;     //96pi/512
  assign cos2[96]  =  7'b0011100;     //96pi/512
  assign sin2[97]  =  7'b1110001;     //97pi/512
  assign cos2[97]  =  7'b0011100;     //97pi/512
  assign sin2[98]  =  7'b1110001;     //98pi/512
  assign cos2[98]  =  7'b0011100;     //98pi/512
  assign sin2[99]  =  7'b1110001;     //99pi/512
  assign cos2[99]  =  7'b0011100;     //99pi/512
  assign sin2[100]  =  7'b1110001;     //100pi/512
  assign cos2[100]  =  7'b0011100;     //100pi/512
  assign sin2[101]  =  7'b1110001;     //101pi/512
  assign cos2[101]  =  7'b0011100;     //101pi/512
  assign sin2[102]  =  7'b1110001;     //102pi/512
  assign cos2[102]  =  7'b0011100;     //102pi/512
  assign sin2[103]  =  7'b1110001;     //103pi/512
  assign cos2[103]  =  7'b0011011;     //103pi/512
  assign sin2[104]  =  7'b1110000;     //104pi/512
  assign cos2[104]  =  7'b0011011;     //104pi/512
  assign sin2[105]  =  7'b1110000;     //105pi/512
  assign cos2[105]  =  7'b0011011;     //105pi/512
  assign sin2[106]  =  7'b1110000;     //106pi/512
  assign cos2[106]  =  7'b0011011;     //106pi/512
  assign sin2[107]  =  7'b1110000;     //107pi/512
  assign cos2[107]  =  7'b0011011;     //107pi/512
  assign sin2[108]  =  7'b1110000;     //108pi/512
  assign cos2[108]  =  7'b0011011;     //108pi/512
  assign sin2[109]  =  7'b1110000;     //109pi/512
  assign cos2[109]  =  7'b0011011;     //109pi/512
  assign sin2[110]  =  7'b1110000;     //110pi/512
  assign cos2[110]  =  7'b0011011;     //110pi/512
  assign sin2[111]  =  7'b1101111;     //111pi/512
  assign cos2[111]  =  7'b0011011;     //111pi/512
  assign sin2[112]  =  7'b1101111;     //112pi/512
  assign cos2[112]  =  7'b0011011;     //112pi/512
  assign sin2[113]  =  7'b1101111;     //113pi/512
  assign cos2[113]  =  7'b0011011;     //113pi/512
  assign sin2[114]  =  7'b1101111;     //114pi/512
  assign cos2[114]  =  7'b0011011;     //114pi/512
  assign sin2[115]  =  7'b1101111;     //115pi/512
  assign cos2[115]  =  7'b0011011;     //115pi/512
  assign sin2[116]  =  7'b1101111;     //116pi/512
  assign cos2[116]  =  7'b0011010;     //116pi/512
  assign sin2[117]  =  7'b1101111;     //117pi/512
  assign cos2[117]  =  7'b0011010;     //117pi/512
  assign sin2[118]  =  7'b1101110;     //118pi/512
  assign cos2[118]  =  7'b0011010;     //118pi/512
  assign sin2[119]  =  7'b1101110;     //119pi/512
  assign cos2[119]  =  7'b0011010;     //119pi/512
  assign sin2[120]  =  7'b1101110;     //120pi/512
  assign cos2[120]  =  7'b0011010;     //120pi/512
  assign sin2[121]  =  7'b1101110;     //121pi/512
  assign cos2[121]  =  7'b0011010;     //121pi/512
  assign sin2[122]  =  7'b1101110;     //122pi/512
  assign cos2[122]  =  7'b0011010;     //122pi/512
  assign sin2[123]  =  7'b1101110;     //123pi/512
  assign cos2[123]  =  7'b0011010;     //123pi/512
  assign sin2[124]  =  7'b1101110;     //124pi/512
  assign cos2[124]  =  7'b0011010;     //124pi/512
  assign sin2[125]  =  7'b1101110;     //125pi/512
  assign cos2[125]  =  7'b0011010;     //125pi/512
  assign sin2[126]  =  7'b1101101;     //126pi/512
  assign cos2[126]  =  7'b0011010;     //126pi/512
  assign sin2[127]  =  7'b1101101;     //127pi/512
  assign cos2[127]  =  7'b0011001;     //127pi/512
  assign sin2[128]  =  7'b1101101;     //128pi/512
  assign cos2[128]  =  7'b0011001;     //128pi/512
  assign sin2[129]  =  7'b1101101;     //129pi/512
  assign cos2[129]  =  7'b0011001;     //129pi/512
  assign sin2[130]  =  7'b1101101;     //130pi/512
  assign cos2[130]  =  7'b0011001;     //130pi/512
  assign sin2[131]  =  7'b1101101;     //131pi/512
  assign cos2[131]  =  7'b0011001;     //131pi/512
  assign sin2[132]  =  7'b1101101;     //132pi/512
  assign cos2[132]  =  7'b0011001;     //132pi/512
  assign sin2[133]  =  7'b1101101;     //133pi/512
  assign cos2[133]  =  7'b0011001;     //133pi/512
  assign sin2[134]  =  7'b1101100;     //134pi/512
  assign cos2[134]  =  7'b0011001;     //134pi/512
  assign sin2[135]  =  7'b1101100;     //135pi/512
  assign cos2[135]  =  7'b0011001;     //135pi/512
  assign sin2[136]  =  7'b1101100;     //136pi/512
  assign cos2[136]  =  7'b0011001;     //136pi/512
  assign sin2[137]  =  7'b1101100;     //137pi/512
  assign cos2[137]  =  7'b0011001;     //137pi/512
  assign sin2[138]  =  7'b1101100;     //138pi/512
  assign cos2[138]  =  7'b0011000;     //138pi/512
  assign sin2[139]  =  7'b1101100;     //139pi/512
  assign cos2[139]  =  7'b0011000;     //139pi/512
  assign sin2[140]  =  7'b1101100;     //140pi/512
  assign cos2[140]  =  7'b0011000;     //140pi/512
  assign sin2[141]  =  7'b1101100;     //141pi/512
  assign cos2[141]  =  7'b0011000;     //141pi/512
  assign sin2[142]  =  7'b1101011;     //142pi/512
  assign cos2[142]  =  7'b0011000;     //142pi/512
  assign sin2[143]  =  7'b1101011;     //143pi/512
  assign cos2[143]  =  7'b0011000;     //143pi/512
  assign sin2[144]  =  7'b1101011;     //144pi/512
  assign cos2[144]  =  7'b0011000;     //144pi/512
  assign sin2[145]  =  7'b1101011;     //145pi/512
  assign cos2[145]  =  7'b0011000;     //145pi/512
  assign sin2[146]  =  7'b1101011;     //146pi/512
  assign cos2[146]  =  7'b0011000;     //146pi/512
  assign sin2[147]  =  7'b1101011;     //147pi/512
  assign cos2[147]  =  7'b0011000;     //147pi/512
  assign sin2[148]  =  7'b1101011;     //148pi/512
  assign cos2[148]  =  7'b0010111;     //148pi/512
  assign sin2[149]  =  7'b1101011;     //149pi/512
  assign cos2[149]  =  7'b0010111;     //149pi/512
  assign sin2[150]  =  7'b1101011;     //150pi/512
  assign cos2[150]  =  7'b0010111;     //150pi/512
  assign sin2[151]  =  7'b1101010;     //151pi/512
  assign cos2[151]  =  7'b0010111;     //151pi/512
  assign sin2[152]  =  7'b1101010;     //152pi/512
  assign cos2[152]  =  7'b0010111;     //152pi/512
  assign sin2[153]  =  7'b1101010;     //153pi/512
  assign cos2[153]  =  7'b0010111;     //153pi/512
  assign sin2[154]  =  7'b1101010;     //154pi/512
  assign cos2[154]  =  7'b0010111;     //154pi/512
  assign sin2[155]  =  7'b1101010;     //155pi/512
  assign cos2[155]  =  7'b0010111;     //155pi/512
  assign sin2[156]  =  7'b1101010;     //156pi/512
  assign cos2[156]  =  7'b0010111;     //156pi/512
  assign sin2[157]  =  7'b1101010;     //157pi/512
  assign cos2[157]  =  7'b0010110;     //157pi/512
  assign sin2[158]  =  7'b1101010;     //158pi/512
  assign cos2[158]  =  7'b0010110;     //158pi/512
  assign sin2[159]  =  7'b1101001;     //159pi/512
  assign cos2[159]  =  7'b0010110;     //159pi/512
  assign sin2[160]  =  7'b1101001;     //160pi/512
  assign cos2[160]  =  7'b0010110;     //160pi/512
  assign sin2[161]  =  7'b1101001;     //161pi/512
  assign cos2[161]  =  7'b0010110;     //161pi/512
  assign sin2[162]  =  7'b1101001;     //162pi/512
  assign cos2[162]  =  7'b0010110;     //162pi/512
  assign sin2[163]  =  7'b1101001;     //163pi/512
  assign cos2[163]  =  7'b0010110;     //163pi/512
  assign sin2[164]  =  7'b1101001;     //164pi/512
  assign cos2[164]  =  7'b0010110;     //164pi/512
  assign sin2[165]  =  7'b1101001;     //165pi/512
  assign cos2[165]  =  7'b0010110;     //165pi/512
  assign sin2[166]  =  7'b1101001;     //166pi/512
  assign cos2[166]  =  7'b0010101;     //166pi/512
  assign sin2[167]  =  7'b1101001;     //167pi/512
  assign cos2[167]  =  7'b0010101;     //167pi/512
  assign sin2[168]  =  7'b1101001;     //168pi/512
  assign cos2[168]  =  7'b0010101;     //168pi/512
  assign sin2[169]  =  7'b1101000;     //169pi/512
  assign cos2[169]  =  7'b0010101;     //169pi/512
  assign sin2[170]  =  7'b1101000;     //170pi/512
  assign cos2[170]  =  7'b0010101;     //170pi/512
  assign sin2[171]  =  7'b1101000;     //171pi/512
  assign cos2[171]  =  7'b0010101;     //171pi/512
  assign sin2[172]  =  7'b1101000;     //172pi/512
  assign cos2[172]  =  7'b0010101;     //172pi/512
  assign sin2[173]  =  7'b1101000;     //173pi/512
  assign cos2[173]  =  7'b0010101;     //173pi/512
  assign sin2[174]  =  7'b1101000;     //174pi/512
  assign cos2[174]  =  7'b0010101;     //174pi/512
  assign sin2[175]  =  7'b1101000;     //175pi/512
  assign cos2[175]  =  7'b0010100;     //175pi/512
  assign sin2[176]  =  7'b1101000;     //176pi/512
  assign cos2[176]  =  7'b0010100;     //176pi/512
  assign sin2[177]  =  7'b1101000;     //177pi/512
  assign cos2[177]  =  7'b0010100;     //177pi/512
  assign sin2[178]  =  7'b1100111;     //178pi/512
  assign cos2[178]  =  7'b0010100;     //178pi/512
  assign sin2[179]  =  7'b1100111;     //179pi/512
  assign cos2[179]  =  7'b0010100;     //179pi/512
  assign sin2[180]  =  7'b1100111;     //180pi/512
  assign cos2[180]  =  7'b0010100;     //180pi/512
  assign sin2[181]  =  7'b1100111;     //181pi/512
  assign cos2[181]  =  7'b0010100;     //181pi/512
  assign sin2[182]  =  7'b1100111;     //182pi/512
  assign cos2[182]  =  7'b0010100;     //182pi/512
  assign sin2[183]  =  7'b1100111;     //183pi/512
  assign cos2[183]  =  7'b0010011;     //183pi/512
  assign sin2[184]  =  7'b1100111;     //184pi/512
  assign cos2[184]  =  7'b0010011;     //184pi/512
  assign sin2[185]  =  7'b1100111;     //185pi/512
  assign cos2[185]  =  7'b0010011;     //185pi/512
  assign sin2[186]  =  7'b1100111;     //186pi/512
  assign cos2[186]  =  7'b0010011;     //186pi/512
  assign sin2[187]  =  7'b1100111;     //187pi/512
  assign cos2[187]  =  7'b0010011;     //187pi/512
  assign sin2[188]  =  7'b1100110;     //188pi/512
  assign cos2[188]  =  7'b0010011;     //188pi/512
  assign sin2[189]  =  7'b1100110;     //189pi/512
  assign cos2[189]  =  7'b0010011;     //189pi/512
  assign sin2[190]  =  7'b1100110;     //190pi/512
  assign cos2[190]  =  7'b0010011;     //190pi/512
  assign sin2[191]  =  7'b1100110;     //191pi/512
  assign cos2[191]  =  7'b0010010;     //191pi/512
  assign sin2[192]  =  7'b1100110;     //192pi/512
  assign cos2[192]  =  7'b0010010;     //192pi/512
  assign sin2[193]  =  7'b1100110;     //193pi/512
  assign cos2[193]  =  7'b0010010;     //193pi/512
  assign sin2[194]  =  7'b1100110;     //194pi/512
  assign cos2[194]  =  7'b0010010;     //194pi/512
  assign sin2[195]  =  7'b1100110;     //195pi/512
  assign cos2[195]  =  7'b0010010;     //195pi/512
  assign sin2[196]  =  7'b1100110;     //196pi/512
  assign cos2[196]  =  7'b0010010;     //196pi/512
  assign sin2[197]  =  7'b1100110;     //197pi/512
  assign cos2[197]  =  7'b0010010;     //197pi/512
  assign sin2[198]  =  7'b1100110;     //198pi/512
  assign cos2[198]  =  7'b0010010;     //198pi/512
  assign sin2[199]  =  7'b1100101;     //199pi/512
  assign cos2[199]  =  7'b0010001;     //199pi/512
  assign sin2[200]  =  7'b1100101;     //200pi/512
  assign cos2[200]  =  7'b0010001;     //200pi/512
  assign sin2[201]  =  7'b1100101;     //201pi/512
  assign cos2[201]  =  7'b0010001;     //201pi/512
  assign sin2[202]  =  7'b1100101;     //202pi/512
  assign cos2[202]  =  7'b0010001;     //202pi/512
  assign sin2[203]  =  7'b1100101;     //203pi/512
  assign cos2[203]  =  7'b0010001;     //203pi/512
  assign sin2[204]  =  7'b1100101;     //204pi/512
  assign cos2[204]  =  7'b0010001;     //204pi/512
  assign sin2[205]  =  7'b1100101;     //205pi/512
  assign cos2[205]  =  7'b0010001;     //205pi/512
  assign sin2[206]  =  7'b1100101;     //206pi/512
  assign cos2[206]  =  7'b0010000;     //206pi/512
  assign sin2[207]  =  7'b1100101;     //207pi/512
  assign cos2[207]  =  7'b0010000;     //207pi/512
  assign sin2[208]  =  7'b1100101;     //208pi/512
  assign cos2[208]  =  7'b0010000;     //208pi/512
  assign sin2[209]  =  7'b1100101;     //209pi/512
  assign cos2[209]  =  7'b0010000;     //209pi/512
  assign sin2[210]  =  7'b1100101;     //210pi/512
  assign cos2[210]  =  7'b0010000;     //210pi/512
  assign sin2[211]  =  7'b1100100;     //211pi/512
  assign cos2[211]  =  7'b0010000;     //211pi/512
  assign sin2[212]  =  7'b1100100;     //212pi/512
  assign cos2[212]  =  7'b0010000;     //212pi/512
  assign sin2[213]  =  7'b1100100;     //213pi/512
  assign cos2[213]  =  7'b0010000;     //213pi/512
  assign sin2[214]  =  7'b1100100;     //214pi/512
  assign cos2[214]  =  7'b0001111;     //214pi/512
  assign sin2[215]  =  7'b1100100;     //215pi/512
  assign cos2[215]  =  7'b0001111;     //215pi/512
  assign sin2[216]  =  7'b1100100;     //216pi/512
  assign cos2[216]  =  7'b0001111;     //216pi/512
  assign sin2[217]  =  7'b1100100;     //217pi/512
  assign cos2[217]  =  7'b0001111;     //217pi/512
  assign sin2[218]  =  7'b1100100;     //218pi/512
  assign cos2[218]  =  7'b0001111;     //218pi/512
  assign sin2[219]  =  7'b1100100;     //219pi/512
  assign cos2[219]  =  7'b0001111;     //219pi/512
  assign sin2[220]  =  7'b1100100;     //220pi/512
  assign cos2[220]  =  7'b0001111;     //220pi/512
  assign sin2[221]  =  7'b1100100;     //221pi/512
  assign cos2[221]  =  7'b0001110;     //221pi/512
  assign sin2[222]  =  7'b1100100;     //222pi/512
  assign cos2[222]  =  7'b0001110;     //222pi/512
  assign sin2[223]  =  7'b1100100;     //223pi/512
  assign cos2[223]  =  7'b0001110;     //223pi/512
  assign sin2[224]  =  7'b1100011;     //224pi/512
  assign cos2[224]  =  7'b0001110;     //224pi/512
  assign sin2[225]  =  7'b1100011;     //225pi/512
  assign cos2[225]  =  7'b0001110;     //225pi/512
  assign sin2[226]  =  7'b1100011;     //226pi/512
  assign cos2[226]  =  7'b0001110;     //226pi/512
  assign sin2[227]  =  7'b1100011;     //227pi/512
  assign cos2[227]  =  7'b0001110;     //227pi/512
  assign sin2[228]  =  7'b1100011;     //228pi/512
  assign cos2[228]  =  7'b0001101;     //228pi/512
  assign sin2[229]  =  7'b1100011;     //229pi/512
  assign cos2[229]  =  7'b0001101;     //229pi/512
  assign sin2[230]  =  7'b1100011;     //230pi/512
  assign cos2[230]  =  7'b0001101;     //230pi/512
  assign sin2[231]  =  7'b1100011;     //231pi/512
  assign cos2[231]  =  7'b0001101;     //231pi/512
  assign sin2[232]  =  7'b1100011;     //232pi/512
  assign cos2[232]  =  7'b0001101;     //232pi/512
  assign sin2[233]  =  7'b1100011;     //233pi/512
  assign cos2[233]  =  7'b0001101;     //233pi/512
  assign sin2[234]  =  7'b1100011;     //234pi/512
  assign cos2[234]  =  7'b0001101;     //234pi/512
  assign sin2[235]  =  7'b1100011;     //235pi/512
  assign cos2[235]  =  7'b0001100;     //235pi/512
  assign sin2[236]  =  7'b1100011;     //236pi/512
  assign cos2[236]  =  7'b0001100;     //236pi/512
  assign sin2[237]  =  7'b1100011;     //237pi/512
  assign cos2[237]  =  7'b0001100;     //237pi/512
  assign sin2[238]  =  7'b1100011;     //238pi/512
  assign cos2[238]  =  7'b0001100;     //238pi/512
  assign sin2[239]  =  7'b1100010;     //239pi/512
  assign cos2[239]  =  7'b0001100;     //239pi/512
  assign sin2[240]  =  7'b1100010;     //240pi/512
  assign cos2[240]  =  7'b0001100;     //240pi/512
  assign sin2[241]  =  7'b1100010;     //241pi/512
  assign cos2[241]  =  7'b0001100;     //241pi/512
  assign sin2[242]  =  7'b1100010;     //242pi/512
  assign cos2[242]  =  7'b0001011;     //242pi/512
  assign sin2[243]  =  7'b1100010;     //243pi/512
  assign cos2[243]  =  7'b0001011;     //243pi/512
  assign sin2[244]  =  7'b1100010;     //244pi/512
  assign cos2[244]  =  7'b0001011;     //244pi/512
  assign sin2[245]  =  7'b1100010;     //245pi/512
  assign cos2[245]  =  7'b0001011;     //245pi/512
  assign sin2[246]  =  7'b1100010;     //246pi/512
  assign cos2[246]  =  7'b0001011;     //246pi/512
  assign sin2[247]  =  7'b1100010;     //247pi/512
  assign cos2[247]  =  7'b0001011;     //247pi/512
  assign sin2[248]  =  7'b1100010;     //248pi/512
  assign cos2[248]  =  7'b0001011;     //248pi/512
  assign sin2[249]  =  7'b1100010;     //249pi/512
  assign cos2[249]  =  7'b0001010;     //249pi/512
  assign sin2[250]  =  7'b1100010;     //250pi/512
  assign cos2[250]  =  7'b0001010;     //250pi/512
  assign sin2[251]  =  7'b1100010;     //251pi/512
  assign cos2[251]  =  7'b0001010;     //251pi/512
  assign sin2[252]  =  7'b1100010;     //252pi/512
  assign cos2[252]  =  7'b0001010;     //252pi/512
  assign sin2[253]  =  7'b1100010;     //253pi/512
  assign cos2[253]  =  7'b0001010;     //253pi/512
  assign sin2[254]  =  7'b1100010;     //254pi/512
  assign cos2[254]  =  7'b0001010;     //254pi/512
  assign sin2[255]  =  7'b1100010;     //255pi/512
  assign cos2[255]  =  7'b0001010;     //255pi/512
  assign sin2[256]  =  7'b1100010;     //256pi/512
  assign cos2[256]  =  7'b0001001;     //256pi/512
  assign sin2[257]  =  7'b1100010;     //257pi/512
  assign cos2[257]  =  7'b0001001;     //257pi/512
  assign sin2[258]  =  7'b1100001;     //258pi/512
  assign cos2[258]  =  7'b0001001;     //258pi/512
  assign sin2[259]  =  7'b1100001;     //259pi/512
  assign cos2[259]  =  7'b0001001;     //259pi/512
  assign sin2[260]  =  7'b1100001;     //260pi/512
  assign cos2[260]  =  7'b0001001;     //260pi/512
  assign sin2[261]  =  7'b1100001;     //261pi/512
  assign cos2[261]  =  7'b0001001;     //261pi/512
  assign sin2[262]  =  7'b1100001;     //262pi/512
  assign cos2[262]  =  7'b0001000;     //262pi/512
  assign sin2[263]  =  7'b1100001;     //263pi/512
  assign cos2[263]  =  7'b0001000;     //263pi/512
  assign sin2[264]  =  7'b1100001;     //264pi/512
  assign cos2[264]  =  7'b0001000;     //264pi/512
  assign sin2[265]  =  7'b1100001;     //265pi/512
  assign cos2[265]  =  7'b0001000;     //265pi/512
  assign sin2[266]  =  7'b1100001;     //266pi/512
  assign cos2[266]  =  7'b0001000;     //266pi/512
  assign sin2[267]  =  7'b1100001;     //267pi/512
  assign cos2[267]  =  7'b0001000;     //267pi/512
  assign sin2[268]  =  7'b1100001;     //268pi/512
  assign cos2[268]  =  7'b0001000;     //268pi/512
  assign sin2[269]  =  7'b1100001;     //269pi/512
  assign cos2[269]  =  7'b0000111;     //269pi/512
  assign sin2[270]  =  7'b1100001;     //270pi/512
  assign cos2[270]  =  7'b0000111;     //270pi/512
  assign sin2[271]  =  7'b1100001;     //271pi/512
  assign cos2[271]  =  7'b0000111;     //271pi/512
  assign sin2[272]  =  7'b1100001;     //272pi/512
  assign cos2[272]  =  7'b0000111;     //272pi/512
  assign sin2[273]  =  7'b1100001;     //273pi/512
  assign cos2[273]  =  7'b0000111;     //273pi/512
  assign sin2[274]  =  7'b1100001;     //274pi/512
  assign cos2[274]  =  7'b0000111;     //274pi/512
  assign sin2[275]  =  7'b1100001;     //275pi/512
  assign cos2[275]  =  7'b0000111;     //275pi/512
  assign sin2[276]  =  7'b1100001;     //276pi/512
  assign cos2[276]  =  7'b0000110;     //276pi/512
  assign sin2[277]  =  7'b1100001;     //277pi/512
  assign cos2[277]  =  7'b0000110;     //277pi/512
  assign sin2[278]  =  7'b1100001;     //278pi/512
  assign cos2[278]  =  7'b0000110;     //278pi/512
  assign sin2[279]  =  7'b1100001;     //279pi/512
  assign cos2[279]  =  7'b0000110;     //279pi/512
  assign sin2[280]  =  7'b1100001;     //280pi/512
  assign cos2[280]  =  7'b0000110;     //280pi/512
  assign sin2[281]  =  7'b1100001;     //281pi/512
  assign cos2[281]  =  7'b0000110;     //281pi/512
  assign sin2[282]  =  7'b1100001;     //282pi/512
  assign cos2[282]  =  7'b0000101;     //282pi/512
  assign sin2[283]  =  7'b1100001;     //283pi/512
  assign cos2[283]  =  7'b0000101;     //283pi/512
  assign sin2[284]  =  7'b1100000;     //284pi/512
  assign cos2[284]  =  7'b0000101;     //284pi/512
  assign sin2[285]  =  7'b1100000;     //285pi/512
  assign cos2[285]  =  7'b0000101;     //285pi/512
  assign sin2[286]  =  7'b1100000;     //286pi/512
  assign cos2[286]  =  7'b0000101;     //286pi/512
  assign sin2[287]  =  7'b1100000;     //287pi/512
  assign cos2[287]  =  7'b0000101;     //287pi/512
  assign sin2[288]  =  7'b1100000;     //288pi/512
  assign cos2[288]  =  7'b0000101;     //288pi/512
  assign sin2[289]  =  7'b1100000;     //289pi/512
  assign cos2[289]  =  7'b0000100;     //289pi/512
  assign sin2[290]  =  7'b1100000;     //290pi/512
  assign cos2[290]  =  7'b0000100;     //290pi/512
  assign sin2[291]  =  7'b1100000;     //291pi/512
  assign cos2[291]  =  7'b0000100;     //291pi/512
  assign sin2[292]  =  7'b1100000;     //292pi/512
  assign cos2[292]  =  7'b0000100;     //292pi/512
  assign sin2[293]  =  7'b1100000;     //293pi/512
  assign cos2[293]  =  7'b0000100;     //293pi/512
  assign sin2[294]  =  7'b1100000;     //294pi/512
  assign cos2[294]  =  7'b0000100;     //294pi/512
  assign sin2[295]  =  7'b1100000;     //295pi/512
  assign cos2[295]  =  7'b0000011;     //295pi/512
  assign sin2[296]  =  7'b1100000;     //296pi/512
  assign cos2[296]  =  7'b0000011;     //296pi/512
  assign sin2[297]  =  7'b1100000;     //297pi/512
  assign cos2[297]  =  7'b0000011;     //297pi/512
  assign sin2[298]  =  7'b1100000;     //298pi/512
  assign cos2[298]  =  7'b0000011;     //298pi/512
  assign sin2[299]  =  7'b1100000;     //299pi/512
  assign cos2[299]  =  7'b0000011;     //299pi/512
  assign sin2[300]  =  7'b1100000;     //300pi/512
  assign cos2[300]  =  7'b0000011;     //300pi/512
  assign sin2[301]  =  7'b1100000;     //301pi/512
  assign cos2[301]  =  7'b0000010;     //301pi/512
  assign sin2[302]  =  7'b1100000;     //302pi/512
  assign cos2[302]  =  7'b0000010;     //302pi/512
  assign sin2[303]  =  7'b1100000;     //303pi/512
  assign cos2[303]  =  7'b0000010;     //303pi/512
  assign sin2[304]  =  7'b1100000;     //304pi/512
  assign cos2[304]  =  7'b0000010;     //304pi/512
  assign sin2[305]  =  7'b1100000;     //305pi/512
  assign cos2[305]  =  7'b0000010;     //305pi/512
  assign sin2[306]  =  7'b1100000;     //306pi/512
  assign cos2[306]  =  7'b0000010;     //306pi/512
  assign sin2[307]  =  7'b1100000;     //307pi/512
  assign cos2[307]  =  7'b0000010;     //307pi/512
  assign sin2[308]  =  7'b1100000;     //308pi/512
  assign cos2[308]  =  7'b0000001;     //308pi/512
  assign sin2[309]  =  7'b1100000;     //309pi/512
  assign cos2[309]  =  7'b0000001;     //309pi/512
  assign sin2[310]  =  7'b1100000;     //310pi/512
  assign cos2[310]  =  7'b0000001;     //310pi/512
  assign sin2[311]  =  7'b1100000;     //311pi/512
  assign cos2[311]  =  7'b0000001;     //311pi/512
  assign sin2[312]  =  7'b1100000;     //312pi/512
  assign cos2[312]  =  7'b0000001;     //312pi/512
  assign sin2[313]  =  7'b1100000;     //313pi/512
  assign cos2[313]  =  7'b0000001;     //313pi/512
  assign sin2[314]  =  7'b1100000;     //314pi/512
  assign cos2[314]  =  7'b0000000;     //314pi/512
  assign sin2[315]  =  7'b1100000;     //315pi/512
  assign cos2[315]  =  7'b0000000;     //315pi/512
  assign sin2[316]  =  7'b1100000;     //316pi/512
  assign cos2[316]  =  7'b0000000;     //316pi/512
  assign sin2[317]  =  7'b1100000;     //317pi/512
  assign cos2[317]  =  7'b0000000;     //317pi/512
  assign sin2[318]  =  7'b1100000;     //318pi/512
  assign cos2[318]  =  7'b0000000;     //318pi/512
  assign sin2[319]  =  7'b1100000;     //319pi/512
  assign cos2[319]  =  7'b0000000;     //319pi/512
  assign sin2[320]  =  7'b1100000;     //320pi/512
  assign cos2[320]  =  7'b0000000;     //320pi/512
  assign sin2[321]  =  7'b1100000;     //321pi/512
  assign cos2[321]  =  7'b0000000;     //321pi/512
  assign sin2[322]  =  7'b1100000;     //322pi/512
  assign cos2[322]  =  7'b0000000;     //322pi/512
  assign sin2[323]  =  7'b1100000;     //323pi/512
  assign cos2[323]  =  7'b0000000;     //323pi/512
  assign sin2[324]  =  7'b1100000;     //324pi/512
  assign cos2[324]  =  7'b1111111;     //324pi/512
  assign sin2[325]  =  7'b1100000;     //325pi/512
  assign cos2[325]  =  7'b1111111;     //325pi/512
  assign sin2[326]  =  7'b1100000;     //326pi/512
  assign cos2[326]  =  7'b1111111;     //326pi/512
  assign sin2[327]  =  7'b1100000;     //327pi/512
  assign cos2[327]  =  7'b1111111;     //327pi/512
  assign sin2[328]  =  7'b1100000;     //328pi/512
  assign cos2[328]  =  7'b1111111;     //328pi/512
  assign sin2[329]  =  7'b1100000;     //329pi/512
  assign cos2[329]  =  7'b1111111;     //329pi/512
  assign sin2[330]  =  7'b1100000;     //330pi/512
  assign cos2[330]  =  7'b1111110;     //330pi/512
  assign sin2[331]  =  7'b1100000;     //331pi/512
  assign cos2[331]  =  7'b1111110;     //331pi/512
  assign sin2[332]  =  7'b1100000;     //332pi/512
  assign cos2[332]  =  7'b1111110;     //332pi/512
  assign sin2[333]  =  7'b1100000;     //333pi/512
  assign cos2[333]  =  7'b1111110;     //333pi/512
  assign sin2[334]  =  7'b1100000;     //334pi/512
  assign cos2[334]  =  7'b1111110;     //334pi/512
  assign sin2[335]  =  7'b1100000;     //335pi/512
  assign cos2[335]  =  7'b1111110;     //335pi/512
  assign sin2[336]  =  7'b1100000;     //336pi/512
  assign cos2[336]  =  7'b1111101;     //336pi/512
  assign sin2[337]  =  7'b1100000;     //337pi/512
  assign cos2[337]  =  7'b1111101;     //337pi/512
  assign sin2[338]  =  7'b1100000;     //338pi/512
  assign cos2[338]  =  7'b1111101;     //338pi/512
  assign sin2[339]  =  7'b1100000;     //339pi/512
  assign cos2[339]  =  7'b1111101;     //339pi/512
  assign sin2[340]  =  7'b1100000;     //340pi/512
  assign cos2[340]  =  7'b1111101;     //340pi/512
  assign sin2[341]  =  7'b1100000;     //341pi/512
  assign cos2[341]  =  7'b1111101;     //341pi/512
  assign sin2[342]  =  7'b1100000;     //342pi/512
  assign cos2[342]  =  7'b1111101;     //342pi/512
  assign sin2[343]  =  7'b1100000;     //343pi/512
  assign cos2[343]  =  7'b1111100;     //343pi/512
  assign sin2[344]  =  7'b1100000;     //344pi/512
  assign cos2[344]  =  7'b1111100;     //344pi/512
  assign sin2[345]  =  7'b1100000;     //345pi/512
  assign cos2[345]  =  7'b1111100;     //345pi/512
  assign sin2[346]  =  7'b1100000;     //346pi/512
  assign cos2[346]  =  7'b1111100;     //346pi/512
  assign sin2[347]  =  7'b1100000;     //347pi/512
  assign cos2[347]  =  7'b1111100;     //347pi/512
  assign sin2[348]  =  7'b1100000;     //348pi/512
  assign cos2[348]  =  7'b1111100;     //348pi/512
  assign sin2[349]  =  7'b1100000;     //349pi/512
  assign cos2[349]  =  7'b1111011;     //349pi/512
  assign sin2[350]  =  7'b1100000;     //350pi/512
  assign cos2[350]  =  7'b1111011;     //350pi/512
  assign sin2[351]  =  7'b1100000;     //351pi/512
  assign cos2[351]  =  7'b1111011;     //351pi/512
  assign sin2[352]  =  7'b1100000;     //352pi/512
  assign cos2[352]  =  7'b1111011;     //352pi/512
  assign sin2[353]  =  7'b1100000;     //353pi/512
  assign cos2[353]  =  7'b1111011;     //353pi/512
  assign sin2[354]  =  7'b1100000;     //354pi/512
  assign cos2[354]  =  7'b1111011;     //354pi/512
  assign sin2[355]  =  7'b1100000;     //355pi/512
  assign cos2[355]  =  7'b1111011;     //355pi/512
  assign sin2[356]  =  7'b1100000;     //356pi/512
  assign cos2[356]  =  7'b1111010;     //356pi/512
  assign sin2[357]  =  7'b1100001;     //357pi/512
  assign cos2[357]  =  7'b1111010;     //357pi/512
  assign sin2[358]  =  7'b1100001;     //358pi/512
  assign cos2[358]  =  7'b1111010;     //358pi/512
  assign sin2[359]  =  7'b1100001;     //359pi/512
  assign cos2[359]  =  7'b1111010;     //359pi/512
  assign sin2[360]  =  7'b1100001;     //360pi/512
  assign cos2[360]  =  7'b1111010;     //360pi/512
  assign sin2[361]  =  7'b1100001;     //361pi/512
  assign cos2[361]  =  7'b1111010;     //361pi/512
  assign sin2[362]  =  7'b1100001;     //362pi/512
  assign cos2[362]  =  7'b1111001;     //362pi/512
  assign sin2[363]  =  7'b1100001;     //363pi/512
  assign cos2[363]  =  7'b1111001;     //363pi/512
  assign sin2[364]  =  7'b1100001;     //364pi/512
  assign cos2[364]  =  7'b1111001;     //364pi/512
  assign sin2[365]  =  7'b1100001;     //365pi/512
  assign cos2[365]  =  7'b1111001;     //365pi/512
  assign sin2[366]  =  7'b1100001;     //366pi/512
  assign cos2[366]  =  7'b1111001;     //366pi/512
  assign sin2[367]  =  7'b1100001;     //367pi/512
  assign cos2[367]  =  7'b1111001;     //367pi/512
  assign sin2[368]  =  7'b1100001;     //368pi/512
  assign cos2[368]  =  7'b1111001;     //368pi/512
  assign sin2[369]  =  7'b1100001;     //369pi/512
  assign cos2[369]  =  7'b1111000;     //369pi/512
  assign sin2[370]  =  7'b1100001;     //370pi/512
  assign cos2[370]  =  7'b1111000;     //370pi/512
  assign sin2[371]  =  7'b1100001;     //371pi/512
  assign cos2[371]  =  7'b1111000;     //371pi/512
  assign sin2[372]  =  7'b1100001;     //372pi/512
  assign cos2[372]  =  7'b1111000;     //372pi/512
  assign sin2[373]  =  7'b1100001;     //373pi/512
  assign cos2[373]  =  7'b1111000;     //373pi/512
  assign sin2[374]  =  7'b1100001;     //374pi/512
  assign cos2[374]  =  7'b1111000;     //374pi/512
  assign sin2[375]  =  7'b1100001;     //375pi/512
  assign cos2[375]  =  7'b1110111;     //375pi/512
  assign sin2[376]  =  7'b1100001;     //376pi/512
  assign cos2[376]  =  7'b1110111;     //376pi/512
  assign sin2[377]  =  7'b1100001;     //377pi/512
  assign cos2[377]  =  7'b1110111;     //377pi/512
  assign sin2[378]  =  7'b1100001;     //378pi/512
  assign cos2[378]  =  7'b1110111;     //378pi/512
  assign sin2[379]  =  7'b1100001;     //379pi/512
  assign cos2[379]  =  7'b1110111;     //379pi/512
  assign sin2[380]  =  7'b1100001;     //380pi/512
  assign cos2[380]  =  7'b1110111;     //380pi/512
  assign sin2[381]  =  7'b1100001;     //381pi/512
  assign cos2[381]  =  7'b1110111;     //381pi/512
  assign sin2[382]  =  7'b1100001;     //382pi/512
  assign cos2[382]  =  7'b1110110;     //382pi/512
  assign sin2[383]  =  7'b1100010;     //383pi/512
  assign cos2[383]  =  7'b1110110;     //383pi/512
  assign sin2[384]  =  7'b1100010;     //384pi/512
  assign cos2[384]  =  7'b1110110;     //384pi/512
  assign sin2[385]  =  7'b1100010;     //385pi/512
  assign cos2[385]  =  7'b1110110;     //385pi/512
  assign sin2[386]  =  7'b1100010;     //386pi/512
  assign cos2[386]  =  7'b1110110;     //386pi/512
  assign sin2[387]  =  7'b1100010;     //387pi/512
  assign cos2[387]  =  7'b1110110;     //387pi/512
  assign sin2[388]  =  7'b1100010;     //388pi/512
  assign cos2[388]  =  7'b1110110;     //388pi/512
  assign sin2[389]  =  7'b1100010;     //389pi/512
  assign cos2[389]  =  7'b1110101;     //389pi/512
  assign sin2[390]  =  7'b1100010;     //390pi/512
  assign cos2[390]  =  7'b1110101;     //390pi/512
  assign sin2[391]  =  7'b1100010;     //391pi/512
  assign cos2[391]  =  7'b1110101;     //391pi/512
  assign sin2[392]  =  7'b1100010;     //392pi/512
  assign cos2[392]  =  7'b1110101;     //392pi/512
  assign sin2[393]  =  7'b1100010;     //393pi/512
  assign cos2[393]  =  7'b1110101;     //393pi/512
  assign sin2[394]  =  7'b1100010;     //394pi/512
  assign cos2[394]  =  7'b1110101;     //394pi/512
  assign sin2[395]  =  7'b1100010;     //395pi/512
  assign cos2[395]  =  7'b1110100;     //395pi/512
  assign sin2[396]  =  7'b1100010;     //396pi/512
  assign cos2[396]  =  7'b1110100;     //396pi/512
  assign sin2[397]  =  7'b1100010;     //397pi/512
  assign cos2[397]  =  7'b1110100;     //397pi/512
  assign sin2[398]  =  7'b1100010;     //398pi/512
  assign cos2[398]  =  7'b1110100;     //398pi/512
  assign sin2[399]  =  7'b1100010;     //399pi/512
  assign cos2[399]  =  7'b1110100;     //399pi/512
  assign sin2[400]  =  7'b1100010;     //400pi/512
  assign cos2[400]  =  7'b1110100;     //400pi/512
  assign sin2[401]  =  7'b1100010;     //401pi/512
  assign cos2[401]  =  7'b1110100;     //401pi/512
  assign sin2[402]  =  7'b1100011;     //402pi/512
  assign cos2[402]  =  7'b1110011;     //402pi/512
  assign sin2[403]  =  7'b1100011;     //403pi/512
  assign cos2[403]  =  7'b1110011;     //403pi/512
  assign sin2[404]  =  7'b1100011;     //404pi/512
  assign cos2[404]  =  7'b1110011;     //404pi/512
  assign sin2[405]  =  7'b1100011;     //405pi/512
  assign cos2[405]  =  7'b1110011;     //405pi/512
  assign sin2[406]  =  7'b1100011;     //406pi/512
  assign cos2[406]  =  7'b1110011;     //406pi/512
  assign sin2[407]  =  7'b1100011;     //407pi/512
  assign cos2[407]  =  7'b1110011;     //407pi/512
  assign sin2[408]  =  7'b1100011;     //408pi/512
  assign cos2[408]  =  7'b1110011;     //408pi/512
  assign sin2[409]  =  7'b1100011;     //409pi/512
  assign cos2[409]  =  7'b1110010;     //409pi/512
  assign sin2[410]  =  7'b1100011;     //410pi/512
  assign cos2[410]  =  7'b1110010;     //410pi/512
  assign sin2[411]  =  7'b1100011;     //411pi/512
  assign cos2[411]  =  7'b1110010;     //411pi/512
  assign sin2[412]  =  7'b1100011;     //412pi/512
  assign cos2[412]  =  7'b1110010;     //412pi/512
  assign sin2[413]  =  7'b1100011;     //413pi/512
  assign cos2[413]  =  7'b1110010;     //413pi/512
  assign sin2[414]  =  7'b1100011;     //414pi/512
  assign cos2[414]  =  7'b1110010;     //414pi/512
  assign sin2[415]  =  7'b1100011;     //415pi/512
  assign cos2[415]  =  7'b1110010;     //415pi/512
  assign sin2[416]  =  7'b1100011;     //416pi/512
  assign cos2[416]  =  7'b1110001;     //416pi/512
  assign sin2[417]  =  7'b1100100;     //417pi/512
  assign cos2[417]  =  7'b1110001;     //417pi/512
  assign sin2[418]  =  7'b1100100;     //418pi/512
  assign cos2[418]  =  7'b1110001;     //418pi/512
  assign sin2[419]  =  7'b1100100;     //419pi/512
  assign cos2[419]  =  7'b1110001;     //419pi/512
  assign sin2[420]  =  7'b1100100;     //420pi/512
  assign cos2[420]  =  7'b1110001;     //420pi/512
  assign sin2[421]  =  7'b1100100;     //421pi/512
  assign cos2[421]  =  7'b1110001;     //421pi/512
  assign sin2[422]  =  7'b1100100;     //422pi/512
  assign cos2[422]  =  7'b1110001;     //422pi/512
  assign sin2[423]  =  7'b1100100;     //423pi/512
  assign cos2[423]  =  7'b1110001;     //423pi/512
  assign sin2[424]  =  7'b1100100;     //424pi/512
  assign cos2[424]  =  7'b1110000;     //424pi/512
  assign sin2[425]  =  7'b1100100;     //425pi/512
  assign cos2[425]  =  7'b1110000;     //425pi/512
  assign sin2[426]  =  7'b1100100;     //426pi/512
  assign cos2[426]  =  7'b1110000;     //426pi/512
  assign sin2[427]  =  7'b1100100;     //427pi/512
  assign cos2[427]  =  7'b1110000;     //427pi/512
  assign sin2[428]  =  7'b1100100;     //428pi/512
  assign cos2[428]  =  7'b1110000;     //428pi/512
  assign sin2[429]  =  7'b1100100;     //429pi/512
  assign cos2[429]  =  7'b1110000;     //429pi/512
  assign sin2[430]  =  7'b1100101;     //430pi/512
  assign cos2[430]  =  7'b1110000;     //430pi/512
  assign sin2[431]  =  7'b1100101;     //431pi/512
  assign cos2[431]  =  7'b1101111;     //431pi/512
  assign sin2[432]  =  7'b1100101;     //432pi/512
  assign cos2[432]  =  7'b1101111;     //432pi/512
  assign sin2[433]  =  7'b1100101;     //433pi/512
  assign cos2[433]  =  7'b1101111;     //433pi/512
  assign sin2[434]  =  7'b1100101;     //434pi/512
  assign cos2[434]  =  7'b1101111;     //434pi/512
  assign sin2[435]  =  7'b1100101;     //435pi/512
  assign cos2[435]  =  7'b1101111;     //435pi/512
  assign sin2[436]  =  7'b1100101;     //436pi/512
  assign cos2[436]  =  7'b1101111;     //436pi/512
  assign sin2[437]  =  7'b1100101;     //437pi/512
  assign cos2[437]  =  7'b1101111;     //437pi/512
  assign sin2[438]  =  7'b1100101;     //438pi/512
  assign cos2[438]  =  7'b1101110;     //438pi/512
  assign sin2[439]  =  7'b1100101;     //439pi/512
  assign cos2[439]  =  7'b1101110;     //439pi/512
  assign sin2[440]  =  7'b1100101;     //440pi/512
  assign cos2[440]  =  7'b1101110;     //440pi/512
  assign sin2[441]  =  7'b1100101;     //441pi/512
  assign cos2[441]  =  7'b1101110;     //441pi/512
  assign sin2[442]  =  7'b1100110;     //442pi/512
  assign cos2[442]  =  7'b1101110;     //442pi/512
  assign sin2[443]  =  7'b1100110;     //443pi/512
  assign cos2[443]  =  7'b1101110;     //443pi/512
  assign sin2[444]  =  7'b1100110;     //444pi/512
  assign cos2[444]  =  7'b1101110;     //444pi/512
  assign sin2[445]  =  7'b1100110;     //445pi/512
  assign cos2[445]  =  7'b1101110;     //445pi/512
  assign sin2[446]  =  7'b1100110;     //446pi/512
  assign cos2[446]  =  7'b1101101;     //446pi/512
  assign sin2[447]  =  7'b1100110;     //447pi/512
  assign cos2[447]  =  7'b1101101;     //447pi/512
  assign sin2[448]  =  7'b1100110;     //448pi/512
  assign cos2[448]  =  7'b1101101;     //448pi/512
  assign sin2[449]  =  7'b1100110;     //449pi/512
  assign cos2[449]  =  7'b1101101;     //449pi/512
  assign sin2[450]  =  7'b1100110;     //450pi/512
  assign cos2[450]  =  7'b1101101;     //450pi/512
  assign sin2[451]  =  7'b1100110;     //451pi/512
  assign cos2[451]  =  7'b1101101;     //451pi/512
  assign sin2[452]  =  7'b1100110;     //452pi/512
  assign cos2[452]  =  7'b1101101;     //452pi/512
  assign sin2[453]  =  7'b1100111;     //453pi/512
  assign cos2[453]  =  7'b1101101;     //453pi/512
  assign sin2[454]  =  7'b1100111;     //454pi/512
  assign cos2[454]  =  7'b1101100;     //454pi/512
  assign sin2[455]  =  7'b1100111;     //455pi/512
  assign cos2[455]  =  7'b1101100;     //455pi/512
  assign sin2[456]  =  7'b1100111;     //456pi/512
  assign cos2[456]  =  7'b1101100;     //456pi/512
  assign sin2[457]  =  7'b1100111;     //457pi/512
  assign cos2[457]  =  7'b1101100;     //457pi/512
  assign sin2[458]  =  7'b1100111;     //458pi/512
  assign cos2[458]  =  7'b1101100;     //458pi/512
  assign sin2[459]  =  7'b1100111;     //459pi/512
  assign cos2[459]  =  7'b1101100;     //459pi/512
  assign sin2[460]  =  7'b1100111;     //460pi/512
  assign cos2[460]  =  7'b1101100;     //460pi/512
  assign sin2[461]  =  7'b1100111;     //461pi/512
  assign cos2[461]  =  7'b1101100;     //461pi/512
  assign sin2[462]  =  7'b1100111;     //462pi/512
  assign cos2[462]  =  7'b1101011;     //462pi/512
  assign sin2[463]  =  7'b1101000;     //463pi/512
  assign cos2[463]  =  7'b1101011;     //463pi/512
  assign sin2[464]  =  7'b1101000;     //464pi/512
  assign cos2[464]  =  7'b1101011;     //464pi/512
  assign sin2[465]  =  7'b1101000;     //465pi/512
  assign cos2[465]  =  7'b1101011;     //465pi/512
  assign sin2[466]  =  7'b1101000;     //466pi/512
  assign cos2[466]  =  7'b1101011;     //466pi/512
  assign sin2[467]  =  7'b1101000;     //467pi/512
  assign cos2[467]  =  7'b1101011;     //467pi/512
  assign sin2[468]  =  7'b1101000;     //468pi/512
  assign cos2[468]  =  7'b1101011;     //468pi/512
  assign sin2[469]  =  7'b1101000;     //469pi/512
  assign cos2[469]  =  7'b1101011;     //469pi/512
  assign sin2[470]  =  7'b1101000;     //470pi/512
  assign cos2[470]  =  7'b1101011;     //470pi/512
  assign sin2[471]  =  7'b1101000;     //471pi/512
  assign cos2[471]  =  7'b1101010;     //471pi/512
  assign sin2[472]  =  7'b1101001;     //472pi/512
  assign cos2[472]  =  7'b1101010;     //472pi/512
  assign sin2[473]  =  7'b1101001;     //473pi/512
  assign cos2[473]  =  7'b1101010;     //473pi/512
  assign sin2[474]  =  7'b1101001;     //474pi/512
  assign cos2[474]  =  7'b1101010;     //474pi/512
  assign sin2[475]  =  7'b1101001;     //475pi/512
  assign cos2[475]  =  7'b1101010;     //475pi/512
  assign sin2[476]  =  7'b1101001;     //476pi/512
  assign cos2[476]  =  7'b1101010;     //476pi/512
  assign sin2[477]  =  7'b1101001;     //477pi/512
  assign cos2[477]  =  7'b1101010;     //477pi/512
  assign sin2[478]  =  7'b1101001;     //478pi/512
  assign cos2[478]  =  7'b1101010;     //478pi/512
  assign sin2[479]  =  7'b1101001;     //479pi/512
  assign cos2[479]  =  7'b1101001;     //479pi/512
  assign sin2[480]  =  7'b1101001;     //480pi/512
  assign cos2[480]  =  7'b1101001;     //480pi/512
  assign sin2[481]  =  7'b1101001;     //481pi/512
  assign cos2[481]  =  7'b1101001;     //481pi/512
  assign sin2[482]  =  7'b1101010;     //482pi/512
  assign cos2[482]  =  7'b1101001;     //482pi/512
  assign sin2[483]  =  7'b1101010;     //483pi/512
  assign cos2[483]  =  7'b1101001;     //483pi/512
  assign sin2[484]  =  7'b1101010;     //484pi/512
  assign cos2[484]  =  7'b1101001;     //484pi/512
  assign sin2[485]  =  7'b1101010;     //485pi/512
  assign cos2[485]  =  7'b1101001;     //485pi/512
  assign sin2[486]  =  7'b1101010;     //486pi/512
  assign cos2[486]  =  7'b1101001;     //486pi/512
  assign sin2[487]  =  7'b1101010;     //487pi/512
  assign cos2[487]  =  7'b1101001;     //487pi/512
  assign sin2[488]  =  7'b1101010;     //488pi/512
  assign cos2[488]  =  7'b1101001;     //488pi/512
  assign sin2[489]  =  7'b1101010;     //489pi/512
  assign cos2[489]  =  7'b1101000;     //489pi/512
  assign sin2[490]  =  7'b1101011;     //490pi/512
  assign cos2[490]  =  7'b1101000;     //490pi/512
  assign sin2[491]  =  7'b1101011;     //491pi/512
  assign cos2[491]  =  7'b1101000;     //491pi/512
  assign sin2[492]  =  7'b1101011;     //492pi/512
  assign cos2[492]  =  7'b1101000;     //492pi/512
  assign sin2[493]  =  7'b1101011;     //493pi/512
  assign cos2[493]  =  7'b1101000;     //493pi/512
  assign sin2[494]  =  7'b1101011;     //494pi/512
  assign cos2[494]  =  7'b1101000;     //494pi/512
  assign sin2[495]  =  7'b1101011;     //495pi/512
  assign cos2[495]  =  7'b1101000;     //495pi/512
  assign sin2[496]  =  7'b1101011;     //496pi/512
  assign cos2[496]  =  7'b1101000;     //496pi/512
  assign sin2[497]  =  7'b1101011;     //497pi/512
  assign cos2[497]  =  7'b1101000;     //497pi/512
  assign sin2[498]  =  7'b1101011;     //498pi/512
  assign cos2[498]  =  7'b1100111;     //498pi/512
  assign sin2[499]  =  7'b1101100;     //499pi/512
  assign cos2[499]  =  7'b1100111;     //499pi/512
  assign sin2[500]  =  7'b1101100;     //500pi/512
  assign cos2[500]  =  7'b1100111;     //500pi/512
  assign sin2[501]  =  7'b1101100;     //501pi/512
  assign cos2[501]  =  7'b1100111;     //501pi/512
  assign sin2[502]  =  7'b1101100;     //502pi/512
  assign cos2[502]  =  7'b1100111;     //502pi/512
  assign sin2[503]  =  7'b1101100;     //503pi/512
  assign cos2[503]  =  7'b1100111;     //503pi/512
  assign sin2[504]  =  7'b1101100;     //504pi/512
  assign cos2[504]  =  7'b1100111;     //504pi/512
  assign sin2[505]  =  7'b1101100;     //505pi/512
  assign cos2[505]  =  7'b1100111;     //505pi/512
  assign sin2[506]  =  7'b1101100;     //506pi/512
  assign cos2[506]  =  7'b1100111;     //506pi/512
  assign sin2[507]  =  7'b1101101;     //507pi/512
  assign cos2[507]  =  7'b1100111;     //507pi/512
  assign sin2[508]  =  7'b1101101;     //508pi/512
  assign cos2[508]  =  7'b1100110;     //508pi/512
  assign sin2[509]  =  7'b1101101;     //509pi/512
  assign cos2[509]  =  7'b1100110;     //509pi/512
  assign sin2[510]  =  7'b1101101;     //510pi/512
  assign cos2[510]  =  7'b1100110;     //510pi/512
  assign sin2[511]  =  7'b1101101;     //511pi/512
  assign cos2[511]  =  7'b1100110;     //511pi/512
endmodule