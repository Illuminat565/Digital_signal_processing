module  TWIDLE_14_bit_STAGE8_1  #(parameter N = 256, SIZE = 8, bit_width_tw = 14) (
    input                               clk,
    input          [SIZE        -2:0]   rd_ptr_angle,
    input                               en, 

    output reg signed [bit_width_tw-1:0]   cos_data,
    output reg signed [bit_width_tw-1:0]   sin_data
 );

reg signed [bit_width_tw-1:0]  cos  [N/2-1:0];
reg signed [bit_width_tw-1:0]  sin  [N/2-1:0];

localparam  coefficient =  $clog2(256/N);

wire [6:0] rd_ptr = rd_ptr_angle << coefficient;

always @(posedge clk) begin
  if (en) begin
    cos_data <= cos [rd_ptr];
    sin_data <= sin [rd_ptr];
  end
end


initial begin
   sin[0]  =  14'b00000000000000;     //0pi/256
   cos[0]  =  14'b01000000000000;     //0pi/256
   sin[1]  =  14'b00010011110001;     //0.1pi/256
   cos[1]  =  14'b00111100110111;     //0.1pi/256
   sin[2]  =  14'b00001010000000;     //0.05pi/256
   cos[2]  =  14'b00111111001101;     //0.05pi/256
   sin[3]  =  14'b00011101000011;     //0.15pi/256
   cos[3]  =  14'b00111001000001;     //0.15pi/256
   sin[4]  =  14'b00000101000001;     //0.025pi/256
   cos[4]  =  14'b00111111110011;     //0.025pi/256
   sin[5]  =  14'b00011000011111;     //0.125pi/256
   cos[5]  =  14'b00111011001000;     //0.125pi/256
   sin[6]  =  14'b00001110111100;     //0.075pi/256
   cos[6]  =  14'b00111110001110;     //0.075pi/256
   sin[7]  =  14'b00100001011100;     //0.175pi/256
   cos[7]  =  14'b00110110100100;     //0.175pi/256
   sin[8]  =  14'b00000010100000;     //0.0125pi/256
   cos[8]  =  14'b00111111111100;     //0.0125pi/256
   sin[9]  =  14'b00010110001001;     //0.1125pi/256
   cos[9]  =  14'b00111100000010;     //0.1125pi/256
   sin[10]  =  14'b00001100011111;     //0.0625pi/256
   cos[10]  =  14'b00111110110001;     //0.0625pi/256
   sin[11]  =  14'b00011111010001;     //0.1625pi/256
   cos[11]  =  14'b00110111110101;     //0.1625pi/256
   sin[12]  =  14'b00000111100001;     //0.0375pi/256
   cos[12]  =  14'b00111111100011;     //0.0375pi/256
   sin[13]  =  14'b00011010110010;     //0.1375pi/256
   cos[13]  =  14'b00111010000111;     //0.1375pi/256
   sin[14]  =  14'b00010001010111;     //0.0875pi/256
   cos[14]  =  14'b00111101100110;     //0.0875pi/256
   sin[15]  =  14'b00100011100011;     //0.1875pi/256
   cos[15]  =  14'b00110101001101;     //0.1875pi/256
   sin[16]  =  14'b00000001010000;     //0.00625pi/256
   cos[16]  =  14'b00111111111111;     //0.00625pi/256
   sin[17]  =  14'b00010100111101;     //0.10625pi/256
   cos[17]  =  14'b00111100011101;     //0.10625pi/256
   sin[18]  =  14'b00001011010000;     //0.05625pi/256
   cos[18]  =  14'b00111111000000;     //0.05625pi/256
   sin[19]  =  14'b00011110001010;     //0.15625pi/256
   cos[19]  =  14'b00111000011100;     //0.15625pi/256
   sin[20]  =  14'b00000110010001;     //0.03125pi/256
   cos[20]  =  14'b00111111101100;     //0.03125pi/256
   sin[21]  =  14'b00011001101001;     //0.13125pi/256
   cos[21]  =  14'b00111010101000;     //0.13125pi/256
   sin[22]  =  14'b00010000001010;     //0.08125pi/256
   cos[22]  =  14'b00111101111011;     //0.08125pi/256
   sin[23]  =  14'b00100010100000;     //0.18125pi/256
   cos[23]  =  14'b00110101111001;     //0.18125pi/256
   sin[24]  =  14'b00000011110001;     //0.01875pi/256
   cos[24]  =  14'b00111111111000;     //0.01875pi/256
   sin[25]  =  14'b00010111010100;     //0.11875pi/256
   cos[25]  =  14'b00111011100110;     //0.11875pi/256
   sin[26]  =  14'b00001101101101;     //0.06875pi/256
   cos[26]  =  14'b00111110100000;     //0.06875pi/256
   sin[27]  =  14'b00100000010111;     //0.16875pi/256
   cos[27]  =  14'b00110111001101;     //0.16875pi/256
   sin[28]  =  14'b00001000110001;     //0.04375pi/256
   cos[28]  =  14'b00111111011001;     //0.04375pi/256
   sin[29]  =  14'b00011011111011;     //0.14375pi/256
   cos[29]  =  14'b00111001100101;     //0.14375pi/256
   sin[30]  =  14'b00010010100101;     //0.09375pi/256
   cos[30]  =  14'b00111101001111;     //0.09375pi/256
   sin[31]  =  14'b00100100100110;     //0.19375pi/256
   cos[31]  =  14'b00110100100000;     //0.19375pi/256
   sin[32]  =  14'b00000000101000;     //0.003125pi/256
   cos[32]  =  14'b00111111111111;     //0.003125pi/256
   sin[33]  =  14'b00010100010111;     //0.10313pi/256
   cos[33]  =  14'b00111100101010;     //0.10313pi/256
   sin[34]  =  14'b00001010101000;     //0.053125pi/256
   cos[34]  =  14'b00111111000111;     //0.053125pi/256
   sin[35]  =  14'b00011101100111;     //0.15313pi/256
   cos[35]  =  14'b00111000101111;     //0.15313pi/256
   sin[36]  =  14'b00000101101001;     //0.028125pi/256
   cos[36]  =  14'b00111111110000;     //0.028125pi/256
   sin[37]  =  14'b00011001000100;     //0.12813pi/256
   cos[37]  =  14'b00111010111000;     //0.12813pi/256
   sin[38]  =  14'b00001111100011;     //0.078125pi/256
   cos[38]  =  14'b00111110000101;     //0.078125pi/256
   sin[39]  =  14'b00100001111110;     //0.17813pi/256
   cos[39]  =  14'b00110110001111;     //0.17813pi/256
   sin[40]  =  14'b00000011001000;     //0.015625pi/256
   cos[40]  =  14'b00111111111011;     //0.015625pi/256
   sin[41]  =  14'b00010110101111;     //0.11563pi/256
   cos[41]  =  14'b00111011110100;     //0.11563pi/256
   sin[42]  =  14'b00001101000110;     //0.065625pi/256
   cos[42]  =  14'b00111110101001;     //0.065625pi/256
   sin[43]  =  14'b00011111110100;     //0.16563pi/256
   cos[43]  =  14'b00110111100001;     //0.16563pi/256
   sin[44]  =  14'b00001000001001;     //0.040625pi/256
   cos[44]  =  14'b00111111011110;     //0.040625pi/256
   sin[45]  =  14'b00011011010111;     //0.14062pi/256
   cos[45]  =  14'b00111001110110;     //0.14062pi/256
   sin[46]  =  14'b00010001111110;     //0.090625pi/256
   cos[46]  =  14'b00111101011011;     //0.090625pi/256
   sin[47]  =  14'b00100100000100;     //0.19063pi/256
   cos[47]  =  14'b00110100110111;     //0.19063pi/256
   sin[48]  =  14'b00000001111000;     //0.009375pi/256
   cos[48]  =  14'b00111111111110;     //0.009375pi/256
   sin[49]  =  14'b00010101100011;     //0.10938pi/256
   cos[49]  =  14'b00111100010000;     //0.10938pi/256
   sin[50]  =  14'b00001011110111;     //0.059375pi/256
   cos[50]  =  14'b00111110111000;     //0.059375pi/256
   sin[51]  =  14'b00011110101110;     //0.15938pi/256
   cos[51]  =  14'b00111000001001;     //0.15938pi/256
   sin[52]  =  14'b00000110111001;     //0.034375pi/256
   cos[52]  =  14'b00111111101000;     //0.034375pi/256
   sin[53]  =  14'b00011010001110;     //0.13437pi/256
   cos[53]  =  14'b00111010011000;     //0.13437pi/256
   sin[54]  =  14'b00010000110001;     //0.084375pi/256
   cos[54]  =  14'b00111101110000;     //0.084375pi/256
   sin[55]  =  14'b00100011000010;     //0.18438pi/256
   cos[55]  =  14'b00110101100011;     //0.18438pi/256
   sin[56]  =  14'b00000100011001;     //0.021875pi/256
   cos[56]  =  14'b00111111110110;     //0.021875pi/256
   sin[57]  =  14'b00010111111010;     //0.12188pi/256
   cos[57]  =  14'b00111011010111;     //0.12188pi/256
   sin[58]  =  14'b00001110010101;     //0.071875pi/256
   cos[58]  =  14'b00111110011000;     //0.071875pi/256
   sin[59]  =  14'b00100000111001;     //0.17188pi/256
   cos[59]  =  14'b00110110111001;     //0.17188pi/256
   sin[60]  =  14'b00001001011001;     //0.046875pi/256
   cos[60]  =  14'b00111111010011;     //0.046875pi/256
   sin[61]  =  14'b00011100011111;     //0.14688pi/256
   cos[61]  =  14'b00111001010011;     //0.14688pi/256
   sin[62]  =  14'b00010011001011;     //0.096875pi/256
   cos[62]  =  14'b00111101000011;     //0.096875pi/256
   sin[63]  =  14'b00100101000110;     //0.19688pi/256
   cos[63]  =  14'b00110100001001;     //0.19688pi/256
   sin[64]  =  14'b00000000010100;     //0.0015625pi/256
   cos[64]  =  14'b00111111111111;     //0.0015625pi/256
   sin[65]  =  14'b00010100000100;     //0.10156pi/256
   cos[65]  =  14'b00111100110001;     //0.10156pi/256
   sin[66]  =  14'b00001010010100;     //0.051563pi/256
   cos[66]  =  14'b00111111001010;     //0.051563pi/256
   sin[67]  =  14'b00011101010101;     //0.15156pi/256
   cos[67]  =  14'b00111000111000;     //0.15156pi/256
   sin[68]  =  14'b00000101010101;     //0.026563pi/256
   cos[68]  =  14'b00111111110001;     //0.026563pi/256
   sin[69]  =  14'b00011000110010;     //0.12656pi/256
   cos[69]  =  14'b00111011000000;     //0.12656pi/256
   sin[70]  =  14'b00001111001111;     //0.076563pi/256
   cos[70]  =  14'b00111110001010;     //0.076563pi/256
   sin[71]  =  14'b00100001101101;     //0.17656pi/256
   cos[71]  =  14'b00110110011001;     //0.17656pi/256
   sin[72]  =  14'b00000010110100;     //0.014063pi/256
   cos[72]  =  14'b00111111111100;     //0.014063pi/256
   sin[73]  =  14'b00010110011100;     //0.11406pi/256
   cos[73]  =  14'b00111011111011;     //0.11406pi/256
   sin[74]  =  14'b00001100110010;     //0.064063pi/256
   cos[74]  =  14'b00111110101101;     //0.064063pi/256
   sin[75]  =  14'b00011111100010;     //0.16406pi/256
   cos[75]  =  14'b00110111101011;     //0.16406pi/256
   sin[76]  =  14'b00000111110101;     //0.039062pi/256
   cos[76]  =  14'b00111111100001;     //0.039062pi/256
   sin[77]  =  14'b00011011000101;     //0.13906pi/256
   cos[77]  =  14'b00111001111111;     //0.13906pi/256
   sin[78]  =  14'b00010001101011;     //0.089063pi/256
   cos[78]  =  14'b00111101100000;     //0.089063pi/256
   sin[79]  =  14'b00100011110100;     //0.18906pi/256
   cos[79]  =  14'b00110101000010;     //0.18906pi/256
   sin[80]  =  14'b00000001100100;     //0.0078125pi/256
   cos[80]  =  14'b00111111111110;     //0.0078125pi/256
   sin[81]  =  14'b00010101010000;     //0.10781pi/256
   cos[81]  =  14'b00111100010111;     //0.10781pi/256
   sin[82]  =  14'b00001011100011;     //0.057813pi/256
   cos[82]  =  14'b00111110111100;     //0.057813pi/256
   sin[83]  =  14'b00011110011100;     //0.15781pi/256
   cos[83]  =  14'b00111000010010;     //0.15781pi/256
   sin[84]  =  14'b00000110100101;     //0.032813pi/256
   cos[84]  =  14'b00111111101010;     //0.032813pi/256
   sin[85]  =  14'b00011001111011;     //0.13281pi/256
   cos[85]  =  14'b00111010100000;     //0.13281pi/256
   sin[86]  =  14'b00010000011101;     //0.082813pi/256
   cos[86]  =  14'b00111101110110;     //0.082813pi/256
   sin[87]  =  14'b00100010110001;     //0.18281pi/256
   cos[87]  =  14'b00110101101110;     //0.18281pi/256
   sin[88]  =  14'b00000100000101;     //0.020313pi/256
   cos[88]  =  14'b00111111110111;     //0.020313pi/256
   sin[89]  =  14'b00010111100111;     //0.12031pi/256
   cos[89]  =  14'b00111011011110;     //0.12031pi/256
   sin[90]  =  14'b00001110000001;     //0.070312pi/256
   cos[90]  =  14'b00111110011100;     //0.070312pi/256
   sin[91]  =  14'b00100000101000;     //0.17031pi/256
   cos[91]  =  14'b00110111000011;     //0.17031pi/256
   sin[92]  =  14'b00001001000101;     //0.045313pi/256
   cos[92]  =  14'b00111111010110;     //0.045313pi/256
   sin[93]  =  14'b00011100001101;     //0.14531pi/256
   cos[93]  =  14'b00111001011100;     //0.14531pi/256
   sin[94]  =  14'b00010010111000;     //0.095313pi/256
   cos[94]  =  14'b00111101001001;     //0.095313pi/256
   sin[95]  =  14'b00100100110110;     //0.19531pi/256
   cos[95]  =  14'b00110100010100;     //0.19531pi/256
   sin[96]  =  14'b00000000111100;     //0.0046875pi/256
   cos[96]  =  14'b00111111111111;     //0.0046875pi/256
   sin[97]  =  14'b00010100101010;     //0.10469pi/256
   cos[97]  =  14'b00111100100100;     //0.10469pi/256
   sin[98]  =  14'b00001010111100;     //0.054688pi/256
   cos[98]  =  14'b00111111000011;     //0.054688pi/256
   sin[99]  =  14'b00011101111001;     //0.15469pi/256
   cos[99]  =  14'b00111000100101;     //0.15469pi/256
   sin[100]  =  14'b00000101111101;     //0.029688pi/256
   cos[100]  =  14'b00111111101110;     //0.029688pi/256
   sin[101]  =  14'b00011001010111;     //0.12969pi/256
   cos[101]  =  14'b00111010110000;     //0.12969pi/256
   sin[102]  =  14'b00001111110110;     //0.079688pi/256
   cos[102]  =  14'b00111110000000;     //0.079688pi/256
   sin[103]  =  14'b00100010001111;     //0.17969pi/256
   cos[103]  =  14'b00110110000100;     //0.17969pi/256
   sin[104]  =  14'b00000011011101;     //0.017188pi/256
   cos[104]  =  14'b00111111111010;     //0.017188pi/256
   sin[105]  =  14'b00010111000010;     //0.11719pi/256
   cos[105]  =  14'b00111011101101;     //0.11719pi/256
   sin[106]  =  14'b00001101011010;     //0.067187pi/256
   cos[106]  =  14'b00111110100101;     //0.067187pi/256
   sin[107]  =  14'b00100000000101;     //0.16719pi/256
   cos[107]  =  14'b00110111010111;     //0.16719pi/256
   sin[108]  =  14'b00001000011101;     //0.042188pi/256
   cos[108]  =  14'b00111111011100;     //0.042188pi/256
   sin[109]  =  14'b00011011101001;     //0.14219pi/256
   cos[109]  =  14'b00111001101110;     //0.14219pi/256
   sin[110]  =  14'b00010010010001;     //0.092188pi/256
   cos[110]  =  14'b00111101010101;     //0.092188pi/256
   sin[111]  =  14'b00100100010101;     //0.19219pi/256
   cos[111]  =  14'b00110100101011;     //0.19219pi/256
   sin[112]  =  14'b00000010001100;     //0.010938pi/256
   cos[112]  =  14'b00111111111101;     //0.010938pi/256
   sin[113]  =  14'b00010101110110;     //0.11094pi/256
   cos[113]  =  14'b00111100001001;     //0.11094pi/256
   sin[114]  =  14'b00001100001011;     //0.060938pi/256
   cos[114]  =  14'b00111110110101;     //0.060938pi/256
   sin[115]  =  14'b00011110111111;     //0.16094pi/256
   cos[115]  =  14'b00110111111111;     //0.16094pi/256
   sin[116]  =  14'b00000111001101;     //0.035938pi/256
   cos[116]  =  14'b00111111100101;     //0.035938pi/256
   sin[117]  =  14'b00011010100000;     //0.13594pi/256
   cos[117]  =  14'b00111010010000;     //0.13594pi/256
   sin[118]  =  14'b00010001000100;     //0.085938pi/256
   cos[118]  =  14'b00111101101011;     //0.085938pi/256
   sin[119]  =  14'b00100011010010;     //0.18594pi/256
   cos[119]  =  14'b00110101011000;     //0.18594pi/256
   sin[120]  =  14'b00000100101101;     //0.023438pi/256
   cos[120]  =  14'b00111111110100;     //0.023438pi/256
   sin[121]  =  14'b00011000001100;     //0.12344pi/256
   cos[121]  =  14'b00111011001111;     //0.12344pi/256
   sin[122]  =  14'b00001110101000;     //0.073438pi/256
   cos[122]  =  14'b00111110010011;     //0.073438pi/256
   sin[123]  =  14'b00100001001010;     //0.17344pi/256
   cos[123]  =  14'b00110110101110;     //0.17344pi/256
   sin[124]  =  14'b00001001101100;     //0.048438pi/256
   cos[124]  =  14'b00111111010000;     //0.048438pi/256
   sin[125]  =  14'b00011100110001;     //0.14844pi/256
   cos[125]  =  14'b00111001001010;     //0.14844pi/256
   sin[126]  =  14'b00010011011110;     //0.098438pi/256
   cos[126]  =  14'b00111100111101;     //0.098438pi/256
   sin[127]  =  14'b00100101010111;     //0.19844pi/256
   cos[127]  =  14'b00110011111101;     //0.19844pi/256
end

endmodule