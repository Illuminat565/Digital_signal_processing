//----------------------------------------------------------------------------
// Example
//----------------------------------------------------------------------------

module mux_2_1
(
  input  [3:0] d0, d1,
  input        sel,
  output [3:0] y
);

  assign y = sel ? d1 : d0;

endmodule

//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module mux_4_1
(
  input  [3:0] d0, d1, d2, d3,
  input  [1:0] sel,
  output [3:0] y
);
   logic [3:0] y1, y2;
   
   mux_2_1 m1 (.d0(d1),.d1(d3),.sel(sel[1]),.y(y1));
   mux_2_1 m2 (.d0(d0),.d1(d2),.sel(sel[1]),.y(y2));
   mux_2_1 m3 (.d0(y2),.d1(y1),.sel(sel[0]),.y(y));


  // Task:
  // Implement mux_4_1 using three instances of mux_2_1


endmodule
