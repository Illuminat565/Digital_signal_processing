module  M_TWIDLE_6_bit #(parameter SIZE =10) (
    input            en_modify, 
    input   [10:0]   rd_ptr_angle,

    output  signed [5:0]   cos_data,
    output  signed [5:0]   sin_data
 );


wire signed [5:0]  cos  [511:0];
wire signed [5:0]  sin  [511:0];

wire signed [5:0]  cos2  [511:0];
wire signed [5:0]  sin2  [511:0];

assign cos_data =   en_modify? cos2 [rd_ptr_angle] : cos [rd_ptr_angle];
assign sin_data =   en_modify? sin2 [rd_ptr_angle] : sin [rd_ptr_angle];

  assign sin[0]  =  6'b000000;     //0pi/512
  assign cos[0]  =  6'b010000;     //0pi/512
  assign sin[1]  =  6'b000000;     //1pi/512
  assign cos[1]  =  6'b001111;     //1pi/512
  assign sin[2]  =  6'b000000;     //2pi/512
  assign cos[2]  =  6'b001111;     //2pi/512
  assign sin[3]  =  6'b000000;     //3pi/512
  assign cos[3]  =  6'b001111;     //3pi/512
  assign sin[4]  =  6'b000000;     //4pi/512
  assign cos[4]  =  6'b001111;     //4pi/512
  assign sin[5]  =  6'b000000;     //5pi/512
  assign cos[5]  =  6'b001111;     //5pi/512
  assign sin[6]  =  6'b111111;     //6pi/512
  assign cos[6]  =  6'b001111;     //6pi/512
  assign sin[7]  =  6'b111111;     //7pi/512
  assign cos[7]  =  6'b001111;     //7pi/512
  assign sin[8]  =  6'b111111;     //8pi/512
  assign cos[8]  =  6'b001111;     //8pi/512
  assign sin[9]  =  6'b111111;     //9pi/512
  assign cos[9]  =  6'b001111;     //9pi/512
  assign sin[10]  =  6'b111111;     //10pi/512
  assign cos[10]  =  6'b001111;     //10pi/512
  assign sin[11]  =  6'b111111;     //11pi/512
  assign cos[11]  =  6'b001111;     //11pi/512
  assign sin[12]  =  6'b111111;     //12pi/512
  assign cos[12]  =  6'b001111;     //12pi/512
  assign sin[13]  =  6'b111111;     //13pi/512
  assign cos[13]  =  6'b001111;     //13pi/512
  assign sin[14]  =  6'b111111;     //14pi/512
  assign cos[14]  =  6'b001111;     //14pi/512
  assign sin[15]  =  6'b111111;     //15pi/512
  assign cos[15]  =  6'b001111;     //15pi/512
  assign sin[16]  =  6'b111110;     //16pi/512
  assign cos[16]  =  6'b001111;     //16pi/512
  assign sin[17]  =  6'b111110;     //17pi/512
  assign cos[17]  =  6'b001111;     //17pi/512
  assign sin[18]  =  6'b111110;     //18pi/512
  assign cos[18]  =  6'b001111;     //18pi/512
  assign sin[19]  =  6'b111110;     //19pi/512
  assign cos[19]  =  6'b001111;     //19pi/512
  assign sin[20]  =  6'b111110;     //20pi/512
  assign cos[20]  =  6'b001111;     //20pi/512
  assign sin[21]  =  6'b111110;     //21pi/512
  assign cos[21]  =  6'b001111;     //21pi/512
  assign sin[22]  =  6'b111110;     //22pi/512
  assign cos[22]  =  6'b001111;     //22pi/512
  assign sin[23]  =  6'b111110;     //23pi/512
  assign cos[23]  =  6'b001111;     //23pi/512
  assign sin[24]  =  6'b111110;     //24pi/512
  assign cos[24]  =  6'b001111;     //24pi/512
  assign sin[25]  =  6'b111110;     //25pi/512
  assign cos[25]  =  6'b001111;     //25pi/512
  assign sin[26]  =  6'b111101;     //26pi/512
  assign cos[26]  =  6'b001111;     //26pi/512
  assign sin[27]  =  6'b111101;     //27pi/512
  assign cos[27]  =  6'b001111;     //27pi/512
  assign sin[28]  =  6'b111101;     //28pi/512
  assign cos[28]  =  6'b001111;     //28pi/512
  assign sin[29]  =  6'b111101;     //29pi/512
  assign cos[29]  =  6'b001111;     //29pi/512
  assign sin[30]  =  6'b111101;     //30pi/512
  assign cos[30]  =  6'b001111;     //30pi/512
  assign sin[31]  =  6'b111101;     //31pi/512
  assign cos[31]  =  6'b001111;     //31pi/512
  assign sin[32]  =  6'b111101;     //32pi/512
  assign cos[32]  =  6'b001111;     //32pi/512
  assign sin[33]  =  6'b111101;     //33pi/512
  assign cos[33]  =  6'b001111;     //33pi/512
  assign sin[34]  =  6'b111101;     //34pi/512
  assign cos[34]  =  6'b001111;     //34pi/512
  assign sin[35]  =  6'b111101;     //35pi/512
  assign cos[35]  =  6'b001111;     //35pi/512
  assign sin[36]  =  6'b111100;     //36pi/512
  assign cos[36]  =  6'b001111;     //36pi/512
  assign sin[37]  =  6'b111100;     //37pi/512
  assign cos[37]  =  6'b001111;     //37pi/512
  assign sin[38]  =  6'b111100;     //38pi/512
  assign cos[38]  =  6'b001111;     //38pi/512
  assign sin[39]  =  6'b111100;     //39pi/512
  assign cos[39]  =  6'b001111;     //39pi/512
  assign sin[40]  =  6'b111100;     //40pi/512
  assign cos[40]  =  6'b001111;     //40pi/512
  assign sin[41]  =  6'b111100;     //41pi/512
  assign cos[41]  =  6'b001111;     //41pi/512
  assign sin[42]  =  6'b111100;     //42pi/512
  assign cos[42]  =  6'b001111;     //42pi/512
  assign sin[43]  =  6'b111100;     //43pi/512
  assign cos[43]  =  6'b001111;     //43pi/512
  assign sin[44]  =  6'b111100;     //44pi/512
  assign cos[44]  =  6'b001111;     //44pi/512
  assign sin[45]  =  6'b111100;     //45pi/512
  assign cos[45]  =  6'b001111;     //45pi/512
  assign sin[46]  =  6'b111100;     //46pi/512
  assign cos[46]  =  6'b001111;     //46pi/512
  assign sin[47]  =  6'b111011;     //47pi/512
  assign cos[47]  =  6'b001111;     //47pi/512
  assign sin[48]  =  6'b111011;     //48pi/512
  assign cos[48]  =  6'b001111;     //48pi/512
  assign sin[49]  =  6'b111011;     //49pi/512
  assign cos[49]  =  6'b001111;     //49pi/512
  assign sin[50]  =  6'b111011;     //50pi/512
  assign cos[50]  =  6'b001111;     //50pi/512
  assign sin[51]  =  6'b111011;     //51pi/512
  assign cos[51]  =  6'b001111;     //51pi/512
  assign sin[52]  =  6'b111011;     //52pi/512
  assign cos[52]  =  6'b001111;     //52pi/512
  assign sin[53]  =  6'b111011;     //53pi/512
  assign cos[53]  =  6'b001111;     //53pi/512
  assign sin[54]  =  6'b111011;     //54pi/512
  assign cos[54]  =  6'b001111;     //54pi/512
  assign sin[55]  =  6'b111011;     //55pi/512
  assign cos[55]  =  6'b001111;     //55pi/512
  assign sin[56]  =  6'b111011;     //56pi/512
  assign cos[56]  =  6'b001111;     //56pi/512
  assign sin[57]  =  6'b111011;     //57pi/512
  assign cos[57]  =  6'b001111;     //57pi/512
  assign sin[58]  =  6'b111010;     //58pi/512
  assign cos[58]  =  6'b001110;     //58pi/512
  assign sin[59]  =  6'b111010;     //59pi/512
  assign cos[59]  =  6'b001110;     //59pi/512
  assign sin[60]  =  6'b111010;     //60pi/512
  assign cos[60]  =  6'b001110;     //60pi/512
  assign sin[61]  =  6'b111010;     //61pi/512
  assign cos[61]  =  6'b001110;     //61pi/512
  assign sin[62]  =  6'b111010;     //62pi/512
  assign cos[62]  =  6'b001110;     //62pi/512
  assign sin[63]  =  6'b111010;     //63pi/512
  assign cos[63]  =  6'b001110;     //63pi/512
  assign sin[64]  =  6'b111010;     //64pi/512
  assign cos[64]  =  6'b001110;     //64pi/512
  assign sin[65]  =  6'b111010;     //65pi/512
  assign cos[65]  =  6'b001110;     //65pi/512
  assign sin[66]  =  6'b111010;     //66pi/512
  assign cos[66]  =  6'b001110;     //66pi/512
  assign sin[67]  =  6'b111010;     //67pi/512
  assign cos[67]  =  6'b001110;     //67pi/512
  assign sin[68]  =  6'b111010;     //68pi/512
  assign cos[68]  =  6'b001110;     //68pi/512
  assign sin[69]  =  6'b111001;     //69pi/512
  assign cos[69]  =  6'b001110;     //69pi/512
  assign sin[70]  =  6'b111001;     //70pi/512
  assign cos[70]  =  6'b001110;     //70pi/512
  assign sin[71]  =  6'b111001;     //71pi/512
  assign cos[71]  =  6'b001110;     //71pi/512
  assign sin[72]  =  6'b111001;     //72pi/512
  assign cos[72]  =  6'b001110;     //72pi/512
  assign sin[73]  =  6'b111001;     //73pi/512
  assign cos[73]  =  6'b001110;     //73pi/512
  assign sin[74]  =  6'b111001;     //74pi/512
  assign cos[74]  =  6'b001110;     //74pi/512
  assign sin[75]  =  6'b111001;     //75pi/512
  assign cos[75]  =  6'b001110;     //75pi/512
  assign sin[76]  =  6'b111001;     //76pi/512
  assign cos[76]  =  6'b001110;     //76pi/512
  assign sin[77]  =  6'b111001;     //77pi/512
  assign cos[77]  =  6'b001110;     //77pi/512
  assign sin[78]  =  6'b111001;     //78pi/512
  assign cos[78]  =  6'b001110;     //78pi/512
  assign sin[79]  =  6'b111001;     //79pi/512
  assign cos[79]  =  6'b001110;     //79pi/512
  assign sin[80]  =  6'b111000;     //80pi/512
  assign cos[80]  =  6'b001110;     //80pi/512
  assign sin[81]  =  6'b111000;     //81pi/512
  assign cos[81]  =  6'b001110;     //81pi/512
  assign sin[82]  =  6'b111000;     //82pi/512
  assign cos[82]  =  6'b001110;     //82pi/512
  assign sin[83]  =  6'b111000;     //83pi/512
  assign cos[83]  =  6'b001101;     //83pi/512
  assign sin[84]  =  6'b111000;     //84pi/512
  assign cos[84]  =  6'b001101;     //84pi/512
  assign sin[85]  =  6'b111000;     //85pi/512
  assign cos[85]  =  6'b001101;     //85pi/512
  assign sin[86]  =  6'b111000;     //86pi/512
  assign cos[86]  =  6'b001101;     //86pi/512
  assign sin[87]  =  6'b111000;     //87pi/512
  assign cos[87]  =  6'b001101;     //87pi/512
  assign sin[88]  =  6'b111000;     //88pi/512
  assign cos[88]  =  6'b001101;     //88pi/512
  assign sin[89]  =  6'b111000;     //89pi/512
  assign cos[89]  =  6'b001101;     //89pi/512
  assign sin[90]  =  6'b111000;     //90pi/512
  assign cos[90]  =  6'b001101;     //90pi/512
  assign sin[91]  =  6'b111000;     //91pi/512
  assign cos[91]  =  6'b001101;     //91pi/512
  assign sin[92]  =  6'b110111;     //92pi/512
  assign cos[92]  =  6'b001101;     //92pi/512
  assign sin[93]  =  6'b110111;     //93pi/512
  assign cos[93]  =  6'b001101;     //93pi/512
  assign sin[94]  =  6'b110111;     //94pi/512
  assign cos[94]  =  6'b001101;     //94pi/512
  assign sin[95]  =  6'b110111;     //95pi/512
  assign cos[95]  =  6'b001101;     //95pi/512
  assign sin[96]  =  6'b110111;     //96pi/512
  assign cos[96]  =  6'b001101;     //96pi/512
  assign sin[97]  =  6'b110111;     //97pi/512
  assign cos[97]  =  6'b001101;     //97pi/512
  assign sin[98]  =  6'b110111;     //98pi/512
  assign cos[98]  =  6'b001101;     //98pi/512
  assign sin[99]  =  6'b110111;     //99pi/512
  assign cos[99]  =  6'b001101;     //99pi/512
  assign sin[100]  =  6'b110111;     //100pi/512
  assign cos[100]  =  6'b001101;     //100pi/512
  assign sin[101]  =  6'b110111;     //101pi/512
  assign cos[101]  =  6'b001101;     //101pi/512
  assign sin[102]  =  6'b110111;     //102pi/512
  assign cos[102]  =  6'b001100;     //102pi/512
  assign sin[103]  =  6'b110111;     //103pi/512
  assign cos[103]  =  6'b001100;     //103pi/512
  assign sin[104]  =  6'b110110;     //104pi/512
  assign cos[104]  =  6'b001100;     //104pi/512
  assign sin[105]  =  6'b110110;     //105pi/512
  assign cos[105]  =  6'b001100;     //105pi/512
  assign sin[106]  =  6'b110110;     //106pi/512
  assign cos[106]  =  6'b001100;     //106pi/512
  assign sin[107]  =  6'b110110;     //107pi/512
  assign cos[107]  =  6'b001100;     //107pi/512
  assign sin[108]  =  6'b110110;     //108pi/512
  assign cos[108]  =  6'b001100;     //108pi/512
  assign sin[109]  =  6'b110110;     //109pi/512
  assign cos[109]  =  6'b001100;     //109pi/512
  assign sin[110]  =  6'b110110;     //110pi/512
  assign cos[110]  =  6'b001100;     //110pi/512
  assign sin[111]  =  6'b110110;     //111pi/512
  assign cos[111]  =  6'b001100;     //111pi/512
  assign sin[112]  =  6'b110110;     //112pi/512
  assign cos[112]  =  6'b001100;     //112pi/512
  assign sin[113]  =  6'b110110;     //113pi/512
  assign cos[113]  =  6'b001100;     //113pi/512
  assign sin[114]  =  6'b110110;     //114pi/512
  assign cos[114]  =  6'b001100;     //114pi/512
  assign sin[115]  =  6'b110110;     //115pi/512
  assign cos[115]  =  6'b001100;     //115pi/512
  assign sin[116]  =  6'b110110;     //116pi/512
  assign cos[116]  =  6'b001100;     //116pi/512
  assign sin[117]  =  6'b110101;     //117pi/512
  assign cos[117]  =  6'b001100;     //117pi/512
  assign sin[118]  =  6'b110101;     //118pi/512
  assign cos[118]  =  6'b001011;     //118pi/512
  assign sin[119]  =  6'b110101;     //119pi/512
  assign cos[119]  =  6'b001011;     //119pi/512
  assign sin[120]  =  6'b110101;     //120pi/512
  assign cos[120]  =  6'b001011;     //120pi/512
  assign sin[121]  =  6'b110101;     //121pi/512
  assign cos[121]  =  6'b001011;     //121pi/512
  assign sin[122]  =  6'b110101;     //122pi/512
  assign cos[122]  =  6'b001011;     //122pi/512
  assign sin[123]  =  6'b110101;     //123pi/512
  assign cos[123]  =  6'b001011;     //123pi/512
  assign sin[124]  =  6'b110101;     //124pi/512
  assign cos[124]  =  6'b001011;     //124pi/512
  assign sin[125]  =  6'b110101;     //125pi/512
  assign cos[125]  =  6'b001011;     //125pi/512
  assign sin[126]  =  6'b110101;     //126pi/512
  assign cos[126]  =  6'b001011;     //126pi/512
  assign sin[127]  =  6'b110101;     //127pi/512
  assign cos[127]  =  6'b001011;     //127pi/512
  assign sin[128]  =  6'b110101;     //128pi/512
  assign cos[128]  =  6'b001011;     //128pi/512
  assign sin[129]  =  6'b110101;     //129pi/512
  assign cos[129]  =  6'b001011;     //129pi/512
  assign sin[130]  =  6'b110101;     //130pi/512
  assign cos[130]  =  6'b001011;     //130pi/512
  assign sin[131]  =  6'b110100;     //131pi/512
  assign cos[131]  =  6'b001011;     //131pi/512
  assign sin[132]  =  6'b110100;     //132pi/512
  assign cos[132]  =  6'b001011;     //132pi/512
  assign sin[133]  =  6'b110100;     //133pi/512
  assign cos[133]  =  6'b001010;     //133pi/512
  assign sin[134]  =  6'b110100;     //134pi/512
  assign cos[134]  =  6'b001010;     //134pi/512
  assign sin[135]  =  6'b110100;     //135pi/512
  assign cos[135]  =  6'b001010;     //135pi/512
  assign sin[136]  =  6'b110100;     //136pi/512
  assign cos[136]  =  6'b001010;     //136pi/512
  assign sin[137]  =  6'b110100;     //137pi/512
  assign cos[137]  =  6'b001010;     //137pi/512
  assign sin[138]  =  6'b110100;     //138pi/512
  assign cos[138]  =  6'b001010;     //138pi/512
  assign sin[139]  =  6'b110100;     //139pi/512
  assign cos[139]  =  6'b001010;     //139pi/512
  assign sin[140]  =  6'b110100;     //140pi/512
  assign cos[140]  =  6'b001010;     //140pi/512
  assign sin[141]  =  6'b110100;     //141pi/512
  assign cos[141]  =  6'b001010;     //141pi/512
  assign sin[142]  =  6'b110100;     //142pi/512
  assign cos[142]  =  6'b001010;     //142pi/512
  assign sin[143]  =  6'b110100;     //143pi/512
  assign cos[143]  =  6'b001010;     //143pi/512
  assign sin[144]  =  6'b110100;     //144pi/512
  assign cos[144]  =  6'b001010;     //144pi/512
  assign sin[145]  =  6'b110100;     //145pi/512
  assign cos[145]  =  6'b001010;     //145pi/512
  assign sin[146]  =  6'b110100;     //146pi/512
  assign cos[146]  =  6'b001001;     //146pi/512
  assign sin[147]  =  6'b110011;     //147pi/512
  assign cos[147]  =  6'b001001;     //147pi/512
  assign sin[148]  =  6'b110011;     //148pi/512
  assign cos[148]  =  6'b001001;     //148pi/512
  assign sin[149]  =  6'b110011;     //149pi/512
  assign cos[149]  =  6'b001001;     //149pi/512
  assign sin[150]  =  6'b110011;     //150pi/512
  assign cos[150]  =  6'b001001;     //150pi/512
  assign sin[151]  =  6'b110011;     //151pi/512
  assign cos[151]  =  6'b001001;     //151pi/512
  assign sin[152]  =  6'b110011;     //152pi/512
  assign cos[152]  =  6'b001001;     //152pi/512
  assign sin[153]  =  6'b110011;     //153pi/512
  assign cos[153]  =  6'b001001;     //153pi/512
  assign sin[154]  =  6'b110011;     //154pi/512
  assign cos[154]  =  6'b001001;     //154pi/512
  assign sin[155]  =  6'b110011;     //155pi/512
  assign cos[155]  =  6'b001001;     //155pi/512
  assign sin[156]  =  6'b110011;     //156pi/512
  assign cos[156]  =  6'b001001;     //156pi/512
  assign sin[157]  =  6'b110011;     //157pi/512
  assign cos[157]  =  6'b001001;     //157pi/512
  assign sin[158]  =  6'b110011;     //158pi/512
  assign cos[158]  =  6'b001001;     //158pi/512
  assign sin[159]  =  6'b110011;     //159pi/512
  assign cos[159]  =  6'b001000;     //159pi/512
  assign sin[160]  =  6'b110011;     //160pi/512
  assign cos[160]  =  6'b001000;     //160pi/512
  assign sin[161]  =  6'b110011;     //161pi/512
  assign cos[161]  =  6'b001000;     //161pi/512
  assign sin[162]  =  6'b110011;     //162pi/512
  assign cos[162]  =  6'b001000;     //162pi/512
  assign sin[163]  =  6'b110011;     //163pi/512
  assign cos[163]  =  6'b001000;     //163pi/512
  assign sin[164]  =  6'b110010;     //164pi/512
  assign cos[164]  =  6'b001000;     //164pi/512
  assign sin[165]  =  6'b110010;     //165pi/512
  assign cos[165]  =  6'b001000;     //165pi/512
  assign sin[166]  =  6'b110010;     //166pi/512
  assign cos[166]  =  6'b001000;     //166pi/512
  assign sin[167]  =  6'b110010;     //167pi/512
  assign cos[167]  =  6'b001000;     //167pi/512
  assign sin[168]  =  6'b110010;     //168pi/512
  assign cos[168]  =  6'b001000;     //168pi/512
  assign sin[169]  =  6'b110010;     //169pi/512
  assign cos[169]  =  6'b001000;     //169pi/512
  assign sin[170]  =  6'b110010;     //170pi/512
  assign cos[170]  =  6'b001000;     //170pi/512
  assign sin[171]  =  6'b110010;     //171pi/512
  assign cos[171]  =  6'b000111;     //171pi/512
  assign sin[172]  =  6'b110010;     //172pi/512
  assign cos[172]  =  6'b000111;     //172pi/512
  assign sin[173]  =  6'b110010;     //173pi/512
  assign cos[173]  =  6'b000111;     //173pi/512
  assign sin[174]  =  6'b110010;     //174pi/512
  assign cos[174]  =  6'b000111;     //174pi/512
  assign sin[175]  =  6'b110010;     //175pi/512
  assign cos[175]  =  6'b000111;     //175pi/512
  assign sin[176]  =  6'b110010;     //176pi/512
  assign cos[176]  =  6'b000111;     //176pi/512
  assign sin[177]  =  6'b110010;     //177pi/512
  assign cos[177]  =  6'b000111;     //177pi/512
  assign sin[178]  =  6'b110010;     //178pi/512
  assign cos[178]  =  6'b000111;     //178pi/512
  assign sin[179]  =  6'b110010;     //179pi/512
  assign cos[179]  =  6'b000111;     //179pi/512
  assign sin[180]  =  6'b110010;     //180pi/512
  assign cos[180]  =  6'b000111;     //180pi/512
  assign sin[181]  =  6'b110010;     //181pi/512
  assign cos[181]  =  6'b000111;     //181pi/512
  assign sin[182]  =  6'b110010;     //182pi/512
  assign cos[182]  =  6'b000111;     //182pi/512
  assign sin[183]  =  6'b110010;     //183pi/512
  assign cos[183]  =  6'b000110;     //183pi/512
  assign sin[184]  =  6'b110010;     //184pi/512
  assign cos[184]  =  6'b000110;     //184pi/512
  assign sin[185]  =  6'b110001;     //185pi/512
  assign cos[185]  =  6'b000110;     //185pi/512
  assign sin[186]  =  6'b110001;     //186pi/512
  assign cos[186]  =  6'b000110;     //186pi/512
  assign sin[187]  =  6'b110001;     //187pi/512
  assign cos[187]  =  6'b000110;     //187pi/512
  assign sin[188]  =  6'b110001;     //188pi/512
  assign cos[188]  =  6'b000110;     //188pi/512
  assign sin[189]  =  6'b110001;     //189pi/512
  assign cos[189]  =  6'b000110;     //189pi/512
  assign sin[190]  =  6'b110001;     //190pi/512
  assign cos[190]  =  6'b000110;     //190pi/512
  assign sin[191]  =  6'b110001;     //191pi/512
  assign cos[191]  =  6'b000110;     //191pi/512
  assign sin[192]  =  6'b110001;     //192pi/512
  assign cos[192]  =  6'b000110;     //192pi/512
  assign sin[193]  =  6'b110001;     //193pi/512
  assign cos[193]  =  6'b000110;     //193pi/512
  assign sin[194]  =  6'b110001;     //194pi/512
  assign cos[194]  =  6'b000101;     //194pi/512
  assign sin[195]  =  6'b110001;     //195pi/512
  assign cos[195]  =  6'b000101;     //195pi/512
  assign sin[196]  =  6'b110001;     //196pi/512
  assign cos[196]  =  6'b000101;     //196pi/512
  assign sin[197]  =  6'b110001;     //197pi/512
  assign cos[197]  =  6'b000101;     //197pi/512
  assign sin[198]  =  6'b110001;     //198pi/512
  assign cos[198]  =  6'b000101;     //198pi/512
  assign sin[199]  =  6'b110001;     //199pi/512
  assign cos[199]  =  6'b000101;     //199pi/512
  assign sin[200]  =  6'b110001;     //200pi/512
  assign cos[200]  =  6'b000101;     //200pi/512
  assign sin[201]  =  6'b110001;     //201pi/512
  assign cos[201]  =  6'b000101;     //201pi/512
  assign sin[202]  =  6'b110001;     //202pi/512
  assign cos[202]  =  6'b000101;     //202pi/512
  assign sin[203]  =  6'b110001;     //203pi/512
  assign cos[203]  =  6'b000101;     //203pi/512
  assign sin[204]  =  6'b110001;     //204pi/512
  assign cos[204]  =  6'b000101;     //204pi/512
  assign sin[205]  =  6'b110001;     //205pi/512
  assign cos[205]  =  6'b000100;     //205pi/512
  assign sin[206]  =  6'b110001;     //206pi/512
  assign cos[206]  =  6'b000100;     //206pi/512
  assign sin[207]  =  6'b110001;     //207pi/512
  assign cos[207]  =  6'b000100;     //207pi/512
  assign sin[208]  =  6'b110001;     //208pi/512
  assign cos[208]  =  6'b000100;     //208pi/512
  assign sin[209]  =  6'b110001;     //209pi/512
  assign cos[209]  =  6'b000100;     //209pi/512
  assign sin[210]  =  6'b110001;     //210pi/512
  assign cos[210]  =  6'b000100;     //210pi/512
  assign sin[211]  =  6'b110001;     //211pi/512
  assign cos[211]  =  6'b000100;     //211pi/512
  assign sin[212]  =  6'b110001;     //212pi/512
  assign cos[212]  =  6'b000100;     //212pi/512
  assign sin[213]  =  6'b110001;     //213pi/512
  assign cos[213]  =  6'b000100;     //213pi/512
  assign sin[214]  =  6'b110001;     //214pi/512
  assign cos[214]  =  6'b000100;     //214pi/512
  assign sin[215]  =  6'b110001;     //215pi/512
  assign cos[215]  =  6'b000011;     //215pi/512
  assign sin[216]  =  6'b110000;     //216pi/512
  assign cos[216]  =  6'b000011;     //216pi/512
  assign sin[217]  =  6'b110000;     //217pi/512
  assign cos[217]  =  6'b000011;     //217pi/512
  assign sin[218]  =  6'b110000;     //218pi/512
  assign cos[218]  =  6'b000011;     //218pi/512
  assign sin[219]  =  6'b110000;     //219pi/512
  assign cos[219]  =  6'b000011;     //219pi/512
  assign sin[220]  =  6'b110000;     //220pi/512
  assign cos[220]  =  6'b000011;     //220pi/512
  assign sin[221]  =  6'b110000;     //221pi/512
  assign cos[221]  =  6'b000011;     //221pi/512
  assign sin[222]  =  6'b110000;     //222pi/512
  assign cos[222]  =  6'b000011;     //222pi/512
  assign sin[223]  =  6'b110000;     //223pi/512
  assign cos[223]  =  6'b000011;     //223pi/512
  assign sin[224]  =  6'b110000;     //224pi/512
  assign cos[224]  =  6'b000011;     //224pi/512
  assign sin[225]  =  6'b110000;     //225pi/512
  assign cos[225]  =  6'b000011;     //225pi/512
  assign sin[226]  =  6'b110000;     //226pi/512
  assign cos[226]  =  6'b000010;     //226pi/512
  assign sin[227]  =  6'b110000;     //227pi/512
  assign cos[227]  =  6'b000010;     //227pi/512
  assign sin[228]  =  6'b110000;     //228pi/512
  assign cos[228]  =  6'b000010;     //228pi/512
  assign sin[229]  =  6'b110000;     //229pi/512
  assign cos[229]  =  6'b000010;     //229pi/512
  assign sin[230]  =  6'b110000;     //230pi/512
  assign cos[230]  =  6'b000010;     //230pi/512
  assign sin[231]  =  6'b110000;     //231pi/512
  assign cos[231]  =  6'b000010;     //231pi/512
  assign sin[232]  =  6'b110000;     //232pi/512
  assign cos[232]  =  6'b000010;     //232pi/512
  assign sin[233]  =  6'b110000;     //233pi/512
  assign cos[233]  =  6'b000010;     //233pi/512
  assign sin[234]  =  6'b110000;     //234pi/512
  assign cos[234]  =  6'b000010;     //234pi/512
  assign sin[235]  =  6'b110000;     //235pi/512
  assign cos[235]  =  6'b000010;     //235pi/512
  assign sin[236]  =  6'b110000;     //236pi/512
  assign cos[236]  =  6'b000001;     //236pi/512
  assign sin[237]  =  6'b110000;     //237pi/512
  assign cos[237]  =  6'b000001;     //237pi/512
  assign sin[238]  =  6'b110000;     //238pi/512
  assign cos[238]  =  6'b000001;     //238pi/512
  assign sin[239]  =  6'b110000;     //239pi/512
  assign cos[239]  =  6'b000001;     //239pi/512
  assign sin[240]  =  6'b110000;     //240pi/512
  assign cos[240]  =  6'b000001;     //240pi/512
  assign sin[241]  =  6'b110000;     //241pi/512
  assign cos[241]  =  6'b000001;     //241pi/512
  assign sin[242]  =  6'b110000;     //242pi/512
  assign cos[242]  =  6'b000001;     //242pi/512
  assign sin[243]  =  6'b110000;     //243pi/512
  assign cos[243]  =  6'b000001;     //243pi/512
  assign sin[244]  =  6'b110000;     //244pi/512
  assign cos[244]  =  6'b000001;     //244pi/512
  assign sin[245]  =  6'b110000;     //245pi/512
  assign cos[245]  =  6'b000001;     //245pi/512
  assign sin[246]  =  6'b110000;     //246pi/512
  assign cos[246]  =  6'b000000;     //246pi/512
  assign sin[247]  =  6'b110000;     //247pi/512
  assign cos[247]  =  6'b000000;     //247pi/512
  assign sin[248]  =  6'b110000;     //248pi/512
  assign cos[248]  =  6'b000000;     //248pi/512
  assign sin[249]  =  6'b110000;     //249pi/512
  assign cos[249]  =  6'b000000;     //249pi/512
  assign sin[250]  =  6'b110000;     //250pi/512
  assign cos[250]  =  6'b000000;     //250pi/512
  assign sin[251]  =  6'b110000;     //251pi/512
  assign cos[251]  =  6'b000000;     //251pi/512
  assign sin[252]  =  6'b110000;     //252pi/512
  assign cos[252]  =  6'b000000;     //252pi/512
  assign sin[253]  =  6'b110000;     //253pi/512
  assign cos[253]  =  6'b000000;     //253pi/512
  assign sin[254]  =  6'b110000;     //254pi/512
  assign cos[254]  =  6'b000000;     //254pi/512
  assign sin[255]  =  6'b110000;     //255pi/512
  assign cos[255]  =  6'b000000;     //255pi/512
  assign sin[256]  =  6'b110000;     //256pi/512
  assign cos[256]  =  6'b000000;     //256pi/512
  assign sin[257]  =  6'b110000;     //257pi/512
  assign cos[257]  =  6'b000000;     //257pi/512
  assign sin[258]  =  6'b110000;     //258pi/512
  assign cos[258]  =  6'b000000;     //258pi/512
  assign sin[259]  =  6'b110000;     //259pi/512
  assign cos[259]  =  6'b000000;     //259pi/512
  assign sin[260]  =  6'b110000;     //260pi/512
  assign cos[260]  =  6'b000000;     //260pi/512
  assign sin[261]  =  6'b110000;     //261pi/512
  assign cos[261]  =  6'b000000;     //261pi/512
  assign sin[262]  =  6'b110000;     //262pi/512
  assign cos[262]  =  6'b111111;     //262pi/512
  assign sin[263]  =  6'b110000;     //263pi/512
  assign cos[263]  =  6'b111111;     //263pi/512
  assign sin[264]  =  6'b110000;     //264pi/512
  assign cos[264]  =  6'b111111;     //264pi/512
  assign sin[265]  =  6'b110000;     //265pi/512
  assign cos[265]  =  6'b111111;     //265pi/512
  assign sin[266]  =  6'b110000;     //266pi/512
  assign cos[266]  =  6'b111111;     //266pi/512
  assign sin[267]  =  6'b110000;     //267pi/512
  assign cos[267]  =  6'b111111;     //267pi/512
  assign sin[268]  =  6'b110000;     //268pi/512
  assign cos[268]  =  6'b111111;     //268pi/512
  assign sin[269]  =  6'b110000;     //269pi/512
  assign cos[269]  =  6'b111111;     //269pi/512
  assign sin[270]  =  6'b110000;     //270pi/512
  assign cos[270]  =  6'b111111;     //270pi/512
  assign sin[271]  =  6'b110000;     //271pi/512
  assign cos[271]  =  6'b111111;     //271pi/512
  assign sin[272]  =  6'b110000;     //272pi/512
  assign cos[272]  =  6'b111110;     //272pi/512
  assign sin[273]  =  6'b110000;     //273pi/512
  assign cos[273]  =  6'b111110;     //273pi/512
  assign sin[274]  =  6'b110000;     //274pi/512
  assign cos[274]  =  6'b111110;     //274pi/512
  assign sin[275]  =  6'b110000;     //275pi/512
  assign cos[275]  =  6'b111110;     //275pi/512
  assign sin[276]  =  6'b110000;     //276pi/512
  assign cos[276]  =  6'b111110;     //276pi/512
  assign sin[277]  =  6'b110000;     //277pi/512
  assign cos[277]  =  6'b111110;     //277pi/512
  assign sin[278]  =  6'b110000;     //278pi/512
  assign cos[278]  =  6'b111110;     //278pi/512
  assign sin[279]  =  6'b110000;     //279pi/512
  assign cos[279]  =  6'b111110;     //279pi/512
  assign sin[280]  =  6'b110000;     //280pi/512
  assign cos[280]  =  6'b111110;     //280pi/512
  assign sin[281]  =  6'b110000;     //281pi/512
  assign cos[281]  =  6'b111110;     //281pi/512
  assign sin[282]  =  6'b110000;     //282pi/512
  assign cos[282]  =  6'b111101;     //282pi/512
  assign sin[283]  =  6'b110000;     //283pi/512
  assign cos[283]  =  6'b111101;     //283pi/512
  assign sin[284]  =  6'b110000;     //284pi/512
  assign cos[284]  =  6'b111101;     //284pi/512
  assign sin[285]  =  6'b110000;     //285pi/512
  assign cos[285]  =  6'b111101;     //285pi/512
  assign sin[286]  =  6'b110000;     //286pi/512
  assign cos[286]  =  6'b111101;     //286pi/512
  assign sin[287]  =  6'b110000;     //287pi/512
  assign cos[287]  =  6'b111101;     //287pi/512
  assign sin[288]  =  6'b110000;     //288pi/512
  assign cos[288]  =  6'b111101;     //288pi/512
  assign sin[289]  =  6'b110000;     //289pi/512
  assign cos[289]  =  6'b111101;     //289pi/512
  assign sin[290]  =  6'b110000;     //290pi/512
  assign cos[290]  =  6'b111101;     //290pi/512
  assign sin[291]  =  6'b110000;     //291pi/512
  assign cos[291]  =  6'b111101;     //291pi/512
  assign sin[292]  =  6'b110000;     //292pi/512
  assign cos[292]  =  6'b111100;     //292pi/512
  assign sin[293]  =  6'b110000;     //293pi/512
  assign cos[293]  =  6'b111100;     //293pi/512
  assign sin[294]  =  6'b110000;     //294pi/512
  assign cos[294]  =  6'b111100;     //294pi/512
  assign sin[295]  =  6'b110000;     //295pi/512
  assign cos[295]  =  6'b111100;     //295pi/512
  assign sin[296]  =  6'b110000;     //296pi/512
  assign cos[296]  =  6'b111100;     //296pi/512
  assign sin[297]  =  6'b110001;     //297pi/512
  assign cos[297]  =  6'b111100;     //297pi/512
  assign sin[298]  =  6'b110001;     //298pi/512
  assign cos[298]  =  6'b111100;     //298pi/512
  assign sin[299]  =  6'b110001;     //299pi/512
  assign cos[299]  =  6'b111100;     //299pi/512
  assign sin[300]  =  6'b110001;     //300pi/512
  assign cos[300]  =  6'b111100;     //300pi/512
  assign sin[301]  =  6'b110001;     //301pi/512
  assign cos[301]  =  6'b111100;     //301pi/512
  assign sin[302]  =  6'b110001;     //302pi/512
  assign cos[302]  =  6'b111100;     //302pi/512
  assign sin[303]  =  6'b110001;     //303pi/512
  assign cos[303]  =  6'b111011;     //303pi/512
  assign sin[304]  =  6'b110001;     //304pi/512
  assign cos[304]  =  6'b111011;     //304pi/512
  assign sin[305]  =  6'b110001;     //305pi/512
  assign cos[305]  =  6'b111011;     //305pi/512
  assign sin[306]  =  6'b110001;     //306pi/512
  assign cos[306]  =  6'b111011;     //306pi/512
  assign sin[307]  =  6'b110001;     //307pi/512
  assign cos[307]  =  6'b111011;     //307pi/512
  assign sin[308]  =  6'b110001;     //308pi/512
  assign cos[308]  =  6'b111011;     //308pi/512
  assign sin[309]  =  6'b110001;     //309pi/512
  assign cos[309]  =  6'b111011;     //309pi/512
  assign sin[310]  =  6'b110001;     //310pi/512
  assign cos[310]  =  6'b111011;     //310pi/512
  assign sin[311]  =  6'b110001;     //311pi/512
  assign cos[311]  =  6'b111011;     //311pi/512
  assign sin[312]  =  6'b110001;     //312pi/512
  assign cos[312]  =  6'b111011;     //312pi/512
  assign sin[313]  =  6'b110001;     //313pi/512
  assign cos[313]  =  6'b111011;     //313pi/512
  assign sin[314]  =  6'b110001;     //314pi/512
  assign cos[314]  =  6'b111010;     //314pi/512
  assign sin[315]  =  6'b110001;     //315pi/512
  assign cos[315]  =  6'b111010;     //315pi/512
  assign sin[316]  =  6'b110001;     //316pi/512
  assign cos[316]  =  6'b111010;     //316pi/512
  assign sin[317]  =  6'b110001;     //317pi/512
  assign cos[317]  =  6'b111010;     //317pi/512
  assign sin[318]  =  6'b110001;     //318pi/512
  assign cos[318]  =  6'b111010;     //318pi/512
  assign sin[319]  =  6'b110001;     //319pi/512
  assign cos[319]  =  6'b111010;     //319pi/512
  assign sin[320]  =  6'b110001;     //320pi/512
  assign cos[320]  =  6'b111010;     //320pi/512
  assign sin[321]  =  6'b110001;     //321pi/512
  assign cos[321]  =  6'b111010;     //321pi/512
  assign sin[322]  =  6'b110001;     //322pi/512
  assign cos[322]  =  6'b111010;     //322pi/512
  assign sin[323]  =  6'b110001;     //323pi/512
  assign cos[323]  =  6'b111010;     //323pi/512
  assign sin[324]  =  6'b110001;     //324pi/512
  assign cos[324]  =  6'b111010;     //324pi/512
  assign sin[325]  =  6'b110001;     //325pi/512
  assign cos[325]  =  6'b111001;     //325pi/512
  assign sin[326]  =  6'b110001;     //326pi/512
  assign cos[326]  =  6'b111001;     //326pi/512
  assign sin[327]  =  6'b110001;     //327pi/512
  assign cos[327]  =  6'b111001;     //327pi/512
  assign sin[328]  =  6'b110010;     //328pi/512
  assign cos[328]  =  6'b111001;     //328pi/512
  assign sin[329]  =  6'b110010;     //329pi/512
  assign cos[329]  =  6'b111001;     //329pi/512
  assign sin[330]  =  6'b110010;     //330pi/512
  assign cos[330]  =  6'b111001;     //330pi/512
  assign sin[331]  =  6'b110010;     //331pi/512
  assign cos[331]  =  6'b111001;     //331pi/512
  assign sin[332]  =  6'b110010;     //332pi/512
  assign cos[332]  =  6'b111001;     //332pi/512
  assign sin[333]  =  6'b110010;     //333pi/512
  assign cos[333]  =  6'b111001;     //333pi/512
  assign sin[334]  =  6'b110010;     //334pi/512
  assign cos[334]  =  6'b111001;     //334pi/512
  assign sin[335]  =  6'b110010;     //335pi/512
  assign cos[335]  =  6'b111001;     //335pi/512
  assign sin[336]  =  6'b110010;     //336pi/512
  assign cos[336]  =  6'b111000;     //336pi/512
  assign sin[337]  =  6'b110010;     //337pi/512
  assign cos[337]  =  6'b111000;     //337pi/512
  assign sin[338]  =  6'b110010;     //338pi/512
  assign cos[338]  =  6'b111000;     //338pi/512
  assign sin[339]  =  6'b110010;     //339pi/512
  assign cos[339]  =  6'b111000;     //339pi/512
  assign sin[340]  =  6'b110010;     //340pi/512
  assign cos[340]  =  6'b111000;     //340pi/512
  assign sin[341]  =  6'b110010;     //341pi/512
  assign cos[341]  =  6'b111000;     //341pi/512
  assign sin[342]  =  6'b110010;     //342pi/512
  assign cos[342]  =  6'b111000;     //342pi/512
  assign sin[343]  =  6'b110010;     //343pi/512
  assign cos[343]  =  6'b111000;     //343pi/512
  assign sin[344]  =  6'b110010;     //344pi/512
  assign cos[344]  =  6'b111000;     //344pi/512
  assign sin[345]  =  6'b110010;     //345pi/512
  assign cos[345]  =  6'b111000;     //345pi/512
  assign sin[346]  =  6'b110010;     //346pi/512
  assign cos[346]  =  6'b111000;     //346pi/512
  assign sin[347]  =  6'b110010;     //347pi/512
  assign cos[347]  =  6'b111000;     //347pi/512
  assign sin[348]  =  6'b110010;     //348pi/512
  assign cos[348]  =  6'b110111;     //348pi/512
  assign sin[349]  =  6'b110011;     //349pi/512
  assign cos[349]  =  6'b110111;     //349pi/512
  assign sin[350]  =  6'b110011;     //350pi/512
  assign cos[350]  =  6'b110111;     //350pi/512
  assign sin[351]  =  6'b110011;     //351pi/512
  assign cos[351]  =  6'b110111;     //351pi/512
  assign sin[352]  =  6'b110011;     //352pi/512
  assign cos[352]  =  6'b110111;     //352pi/512
  assign sin[353]  =  6'b110011;     //353pi/512
  assign cos[353]  =  6'b110111;     //353pi/512
  assign sin[354]  =  6'b110011;     //354pi/512
  assign cos[354]  =  6'b110111;     //354pi/512
  assign sin[355]  =  6'b110011;     //355pi/512
  assign cos[355]  =  6'b110111;     //355pi/512
  assign sin[356]  =  6'b110011;     //356pi/512
  assign cos[356]  =  6'b110111;     //356pi/512
  assign sin[357]  =  6'b110011;     //357pi/512
  assign cos[357]  =  6'b110111;     //357pi/512
  assign sin[358]  =  6'b110011;     //358pi/512
  assign cos[358]  =  6'b110111;     //358pi/512
  assign sin[359]  =  6'b110011;     //359pi/512
  assign cos[359]  =  6'b110111;     //359pi/512
  assign sin[360]  =  6'b110011;     //360pi/512
  assign cos[360]  =  6'b110110;     //360pi/512
  assign sin[361]  =  6'b110011;     //361pi/512
  assign cos[361]  =  6'b110110;     //361pi/512
  assign sin[362]  =  6'b110011;     //362pi/512
  assign cos[362]  =  6'b110110;     //362pi/512
  assign sin[363]  =  6'b110011;     //363pi/512
  assign cos[363]  =  6'b110110;     //363pi/512
  assign sin[364]  =  6'b110011;     //364pi/512
  assign cos[364]  =  6'b110110;     //364pi/512
  assign sin[365]  =  6'b110011;     //365pi/512
  assign cos[365]  =  6'b110110;     //365pi/512
  assign sin[366]  =  6'b110100;     //366pi/512
  assign cos[366]  =  6'b110110;     //366pi/512
  assign sin[367]  =  6'b110100;     //367pi/512
  assign cos[367]  =  6'b110110;     //367pi/512
  assign sin[368]  =  6'b110100;     //368pi/512
  assign cos[368]  =  6'b110110;     //368pi/512
  assign sin[369]  =  6'b110100;     //369pi/512
  assign cos[369]  =  6'b110110;     //369pi/512
  assign sin[370]  =  6'b110100;     //370pi/512
  assign cos[370]  =  6'b110110;     //370pi/512
  assign sin[371]  =  6'b110100;     //371pi/512
  assign cos[371]  =  6'b110110;     //371pi/512
  assign sin[372]  =  6'b110100;     //372pi/512
  assign cos[372]  =  6'b110110;     //372pi/512
  assign sin[373]  =  6'b110100;     //373pi/512
  assign cos[373]  =  6'b110101;     //373pi/512
  assign sin[374]  =  6'b110100;     //374pi/512
  assign cos[374]  =  6'b110101;     //374pi/512
  assign sin[375]  =  6'b110100;     //375pi/512
  assign cos[375]  =  6'b110101;     //375pi/512
  assign sin[376]  =  6'b110100;     //376pi/512
  assign cos[376]  =  6'b110101;     //376pi/512
  assign sin[377]  =  6'b110100;     //377pi/512
  assign cos[377]  =  6'b110101;     //377pi/512
  assign sin[378]  =  6'b110100;     //378pi/512
  assign cos[378]  =  6'b110101;     //378pi/512
  assign sin[379]  =  6'b110100;     //379pi/512
  assign cos[379]  =  6'b110101;     //379pi/512
  assign sin[380]  =  6'b110100;     //380pi/512
  assign cos[380]  =  6'b110101;     //380pi/512
  assign sin[381]  =  6'b110100;     //381pi/512
  assign cos[381]  =  6'b110101;     //381pi/512
  assign sin[382]  =  6'b110101;     //382pi/512
  assign cos[382]  =  6'b110101;     //382pi/512
  assign sin[383]  =  6'b110101;     //383pi/512
  assign cos[383]  =  6'b110101;     //383pi/512
  assign sin[384]  =  6'b110101;     //384pi/512
  assign cos[384]  =  6'b110101;     //384pi/512
  assign sin[385]  =  6'b110101;     //385pi/512
  assign cos[385]  =  6'b110101;     //385pi/512
  assign sin[386]  =  6'b110101;     //386pi/512
  assign cos[386]  =  6'b110101;     //386pi/512
  assign sin[387]  =  6'b110101;     //387pi/512
  assign cos[387]  =  6'b110100;     //387pi/512
  assign sin[388]  =  6'b110101;     //388pi/512
  assign cos[388]  =  6'b110100;     //388pi/512
  assign sin[389]  =  6'b110101;     //389pi/512
  assign cos[389]  =  6'b110100;     //389pi/512
  assign sin[390]  =  6'b110101;     //390pi/512
  assign cos[390]  =  6'b110100;     //390pi/512
  assign sin[391]  =  6'b110101;     //391pi/512
  assign cos[391]  =  6'b110100;     //391pi/512
  assign sin[392]  =  6'b110101;     //392pi/512
  assign cos[392]  =  6'b110100;     //392pi/512
  assign sin[393]  =  6'b110101;     //393pi/512
  assign cos[393]  =  6'b110100;     //393pi/512
  assign sin[394]  =  6'b110101;     //394pi/512
  assign cos[394]  =  6'b110100;     //394pi/512
  assign sin[395]  =  6'b110101;     //395pi/512
  assign cos[395]  =  6'b110100;     //395pi/512
  assign sin[396]  =  6'b110110;     //396pi/512
  assign cos[396]  =  6'b110100;     //396pi/512
  assign sin[397]  =  6'b110110;     //397pi/512
  assign cos[397]  =  6'b110100;     //397pi/512
  assign sin[398]  =  6'b110110;     //398pi/512
  assign cos[398]  =  6'b110100;     //398pi/512
  assign sin[399]  =  6'b110110;     //399pi/512
  assign cos[399]  =  6'b110100;     //399pi/512
  assign sin[400]  =  6'b110110;     //400pi/512
  assign cos[400]  =  6'b110100;     //400pi/512
  assign sin[401]  =  6'b110110;     //401pi/512
  assign cos[401]  =  6'b110100;     //401pi/512
  assign sin[402]  =  6'b110110;     //402pi/512
  assign cos[402]  =  6'b110100;     //402pi/512
  assign sin[403]  =  6'b110110;     //403pi/512
  assign cos[403]  =  6'b110011;     //403pi/512
  assign sin[404]  =  6'b110110;     //404pi/512
  assign cos[404]  =  6'b110011;     //404pi/512
  assign sin[405]  =  6'b110110;     //405pi/512
  assign cos[405]  =  6'b110011;     //405pi/512
  assign sin[406]  =  6'b110110;     //406pi/512
  assign cos[406]  =  6'b110011;     //406pi/512
  assign sin[407]  =  6'b110110;     //407pi/512
  assign cos[407]  =  6'b110011;     //407pi/512
  assign sin[408]  =  6'b110110;     //408pi/512
  assign cos[408]  =  6'b110011;     //408pi/512
  assign sin[409]  =  6'b110111;     //409pi/512
  assign cos[409]  =  6'b110011;     //409pi/512
  assign sin[410]  =  6'b110111;     //410pi/512
  assign cos[410]  =  6'b110011;     //410pi/512
  assign sin[411]  =  6'b110111;     //411pi/512
  assign cos[411]  =  6'b110011;     //411pi/512
  assign sin[412]  =  6'b110111;     //412pi/512
  assign cos[412]  =  6'b110011;     //412pi/512
  assign sin[413]  =  6'b110111;     //413pi/512
  assign cos[413]  =  6'b110011;     //413pi/512
  assign sin[414]  =  6'b110111;     //414pi/512
  assign cos[414]  =  6'b110011;     //414pi/512
  assign sin[415]  =  6'b110111;     //415pi/512
  assign cos[415]  =  6'b110011;     //415pi/512
  assign sin[416]  =  6'b110111;     //416pi/512
  assign cos[416]  =  6'b110011;     //416pi/512
  assign sin[417]  =  6'b110111;     //417pi/512
  assign cos[417]  =  6'b110011;     //417pi/512
  assign sin[418]  =  6'b110111;     //418pi/512
  assign cos[418]  =  6'b110011;     //418pi/512
  assign sin[419]  =  6'b110111;     //419pi/512
  assign cos[419]  =  6'b110011;     //419pi/512
  assign sin[420]  =  6'b110111;     //420pi/512
  assign cos[420]  =  6'b110010;     //420pi/512
  assign sin[421]  =  6'b111000;     //421pi/512
  assign cos[421]  =  6'b110010;     //421pi/512
  assign sin[422]  =  6'b111000;     //422pi/512
  assign cos[422]  =  6'b110010;     //422pi/512
  assign sin[423]  =  6'b111000;     //423pi/512
  assign cos[423]  =  6'b110010;     //423pi/512
  assign sin[424]  =  6'b111000;     //424pi/512
  assign cos[424]  =  6'b110010;     //424pi/512
  assign sin[425]  =  6'b111000;     //425pi/512
  assign cos[425]  =  6'b110010;     //425pi/512
  assign sin[426]  =  6'b111000;     //426pi/512
  assign cos[426]  =  6'b110010;     //426pi/512
  assign sin[427]  =  6'b111000;     //427pi/512
  assign cos[427]  =  6'b110010;     //427pi/512
  assign sin[428]  =  6'b111000;     //428pi/512
  assign cos[428]  =  6'b110010;     //428pi/512
  assign sin[429]  =  6'b111000;     //429pi/512
  assign cos[429]  =  6'b110010;     //429pi/512
  assign sin[430]  =  6'b111000;     //430pi/512
  assign cos[430]  =  6'b110010;     //430pi/512
  assign sin[431]  =  6'b111000;     //431pi/512
  assign cos[431]  =  6'b110010;     //431pi/512
  assign sin[432]  =  6'b111000;     //432pi/512
  assign cos[432]  =  6'b110010;     //432pi/512
  assign sin[433]  =  6'b111001;     //433pi/512
  assign cos[433]  =  6'b110010;     //433pi/512
  assign sin[434]  =  6'b111001;     //434pi/512
  assign cos[434]  =  6'b110010;     //434pi/512
  assign sin[435]  =  6'b111001;     //435pi/512
  assign cos[435]  =  6'b110010;     //435pi/512
  assign sin[436]  =  6'b111001;     //436pi/512
  assign cos[436]  =  6'b110010;     //436pi/512
  assign sin[437]  =  6'b111001;     //437pi/512
  assign cos[437]  =  6'b110010;     //437pi/512
  assign sin[438]  =  6'b111001;     //438pi/512
  assign cos[438]  =  6'b110010;     //438pi/512
  assign sin[439]  =  6'b111001;     //439pi/512
  assign cos[439]  =  6'b110010;     //439pi/512
  assign sin[440]  =  6'b111001;     //440pi/512
  assign cos[440]  =  6'b110010;     //440pi/512
  assign sin[441]  =  6'b111001;     //441pi/512
  assign cos[441]  =  6'b110001;     //441pi/512
  assign sin[442]  =  6'b111001;     //442pi/512
  assign cos[442]  =  6'b110001;     //442pi/512
  assign sin[443]  =  6'b111001;     //443pi/512
  assign cos[443]  =  6'b110001;     //443pi/512
  assign sin[444]  =  6'b111010;     //444pi/512
  assign cos[444]  =  6'b110001;     //444pi/512
  assign sin[445]  =  6'b111010;     //445pi/512
  assign cos[445]  =  6'b110001;     //445pi/512
  assign sin[446]  =  6'b111010;     //446pi/512
  assign cos[446]  =  6'b110001;     //446pi/512
  assign sin[447]  =  6'b111010;     //447pi/512
  assign cos[447]  =  6'b110001;     //447pi/512
  assign sin[448]  =  6'b111010;     //448pi/512
  assign cos[448]  =  6'b110001;     //448pi/512
  assign sin[449]  =  6'b111010;     //449pi/512
  assign cos[449]  =  6'b110001;     //449pi/512
  assign sin[450]  =  6'b111010;     //450pi/512
  assign cos[450]  =  6'b110001;     //450pi/512
  assign sin[451]  =  6'b111010;     //451pi/512
  assign cos[451]  =  6'b110001;     //451pi/512
  assign sin[452]  =  6'b111010;     //452pi/512
  assign cos[452]  =  6'b110001;     //452pi/512
  assign sin[453]  =  6'b111010;     //453pi/512
  assign cos[453]  =  6'b110001;     //453pi/512
  assign sin[454]  =  6'b111010;     //454pi/512
  assign cos[454]  =  6'b110001;     //454pi/512
  assign sin[455]  =  6'b111011;     //455pi/512
  assign cos[455]  =  6'b110001;     //455pi/512
  assign sin[456]  =  6'b111011;     //456pi/512
  assign cos[456]  =  6'b110001;     //456pi/512
  assign sin[457]  =  6'b111011;     //457pi/512
  assign cos[457]  =  6'b110001;     //457pi/512
  assign sin[458]  =  6'b111011;     //458pi/512
  assign cos[458]  =  6'b110001;     //458pi/512
  assign sin[459]  =  6'b111011;     //459pi/512
  assign cos[459]  =  6'b110001;     //459pi/512
  assign sin[460]  =  6'b111011;     //460pi/512
  assign cos[460]  =  6'b110001;     //460pi/512
  assign sin[461]  =  6'b111011;     //461pi/512
  assign cos[461]  =  6'b110001;     //461pi/512
  assign sin[462]  =  6'b111011;     //462pi/512
  assign cos[462]  =  6'b110001;     //462pi/512
  assign sin[463]  =  6'b111011;     //463pi/512
  assign cos[463]  =  6'b110001;     //463pi/512
  assign sin[464]  =  6'b111011;     //464pi/512
  assign cos[464]  =  6'b110001;     //464pi/512
  assign sin[465]  =  6'b111011;     //465pi/512
  assign cos[465]  =  6'b110001;     //465pi/512
  assign sin[466]  =  6'b111100;     //466pi/512
  assign cos[466]  =  6'b110001;     //466pi/512
  assign sin[467]  =  6'b111100;     //467pi/512
  assign cos[467]  =  6'b110001;     //467pi/512
  assign sin[468]  =  6'b111100;     //468pi/512
  assign cos[468]  =  6'b110001;     //468pi/512
  assign sin[469]  =  6'b111100;     //469pi/512
  assign cos[469]  =  6'b110001;     //469pi/512
  assign sin[470]  =  6'b111100;     //470pi/512
  assign cos[470]  =  6'b110001;     //470pi/512
  assign sin[471]  =  6'b111100;     //471pi/512
  assign cos[471]  =  6'b110001;     //471pi/512
  assign sin[472]  =  6'b111100;     //472pi/512
  assign cos[472]  =  6'b110000;     //472pi/512
  assign sin[473]  =  6'b111100;     //473pi/512
  assign cos[473]  =  6'b110000;     //473pi/512
  assign sin[474]  =  6'b111100;     //474pi/512
  assign cos[474]  =  6'b110000;     //474pi/512
  assign sin[475]  =  6'b111100;     //475pi/512
  assign cos[475]  =  6'b110000;     //475pi/512
  assign sin[476]  =  6'b111100;     //476pi/512
  assign cos[476]  =  6'b110000;     //476pi/512
  assign sin[477]  =  6'b111101;     //477pi/512
  assign cos[477]  =  6'b110000;     //477pi/512
  assign sin[478]  =  6'b111101;     //478pi/512
  assign cos[478]  =  6'b110000;     //478pi/512
  assign sin[479]  =  6'b111101;     //479pi/512
  assign cos[479]  =  6'b110000;     //479pi/512
  assign sin[480]  =  6'b111101;     //480pi/512
  assign cos[480]  =  6'b110000;     //480pi/512
  assign sin[481]  =  6'b111101;     //481pi/512
  assign cos[481]  =  6'b110000;     //481pi/512
  assign sin[482]  =  6'b111101;     //482pi/512
  assign cos[482]  =  6'b110000;     //482pi/512
  assign sin[483]  =  6'b111101;     //483pi/512
  assign cos[483]  =  6'b110000;     //483pi/512
  assign sin[484]  =  6'b111101;     //484pi/512
  assign cos[484]  =  6'b110000;     //484pi/512
  assign sin[485]  =  6'b111101;     //485pi/512
  assign cos[485]  =  6'b110000;     //485pi/512
  assign sin[486]  =  6'b111101;     //486pi/512
  assign cos[486]  =  6'b110000;     //486pi/512
  assign sin[487]  =  6'b111110;     //487pi/512
  assign cos[487]  =  6'b110000;     //487pi/512
  assign sin[488]  =  6'b111110;     //488pi/512
  assign cos[488]  =  6'b110000;     //488pi/512
  assign sin[489]  =  6'b111110;     //489pi/512
  assign cos[489]  =  6'b110000;     //489pi/512
  assign sin[490]  =  6'b111110;     //490pi/512
  assign cos[490]  =  6'b110000;     //490pi/512
  assign sin[491]  =  6'b111110;     //491pi/512
  assign cos[491]  =  6'b110000;     //491pi/512
  assign sin[492]  =  6'b111110;     //492pi/512
  assign cos[492]  =  6'b110000;     //492pi/512
  assign sin[493]  =  6'b111110;     //493pi/512
  assign cos[493]  =  6'b110000;     //493pi/512
  assign sin[494]  =  6'b111110;     //494pi/512
  assign cos[494]  =  6'b110000;     //494pi/512
  assign sin[495]  =  6'b111110;     //495pi/512
  assign cos[495]  =  6'b110000;     //495pi/512
  assign sin[496]  =  6'b111110;     //496pi/512
  assign cos[496]  =  6'b110000;     //496pi/512
  assign sin[497]  =  6'b111111;     //497pi/512
  assign cos[497]  =  6'b110000;     //497pi/512
  assign sin[498]  =  6'b111111;     //498pi/512
  assign cos[498]  =  6'b110000;     //498pi/512
  assign sin[499]  =  6'b111111;     //499pi/512
  assign cos[499]  =  6'b110000;     //499pi/512
  assign sin[500]  =  6'b111111;     //500pi/512
  assign cos[500]  =  6'b110000;     //500pi/512
  assign sin[501]  =  6'b111111;     //501pi/512
  assign cos[501]  =  6'b110000;     //501pi/512
  assign sin[502]  =  6'b111111;     //502pi/512
  assign cos[502]  =  6'b110000;     //502pi/512
  assign sin[503]  =  6'b111111;     //503pi/512
  assign cos[503]  =  6'b110000;     //503pi/512
  assign sin[504]  =  6'b111111;     //504pi/512
  assign cos[504]  =  6'b110000;     //504pi/512
  assign sin[505]  =  6'b111111;     //505pi/512
  assign cos[505]  =  6'b110000;     //505pi/512
  assign sin[506]  =  6'b111111;     //506pi/512
  assign cos[506]  =  6'b110000;     //506pi/512
  assign sin[507]  =  6'b000000;     //507pi/512
  assign cos[507]  =  6'b110000;     //507pi/512
  assign sin[508]  =  6'b000000;     //508pi/512
  assign cos[508]  =  6'b110000;     //508pi/512
  assign sin[509]  =  6'b000000;     //509pi/512
  assign cos[509]  =  6'b110000;     //509pi/512
  assign sin[510]  =  6'b000000;     //510pi/512
  assign cos[510]  =  6'b110000;     //510pi/512
  assign sin[511]  =  6'b000000;     //511pi/512
  assign cos[511]  =  6'b110000;     //511pi/512
/////////////////////////////////////////////////////////
  assign sin2[0]  =  6'b000000;     //0pi/512
  assign cos2[0]  =  6'b010000;     //0pi/512
  assign sin2[1]  =  6'b000000;     //1pi/512
  assign cos2[1]  =  6'b001111;     //1pi/512
  assign sin2[2]  =  6'b000000;     //2pi/512
  assign cos2[2]  =  6'b001111;     //2pi/512
  assign sin2[3]  =  6'b000000;     //3pi/512
  assign cos2[3]  =  6'b001111;     //3pi/512
  assign sin2[4]  =  6'b000000;     //4pi/512
  assign cos2[4]  =  6'b001111;     //4pi/512
  assign sin2[5]  =  6'b000000;     //5pi/512
  assign cos2[5]  =  6'b001111;     //5pi/512
  assign sin2[6]  =  6'b000000;     //6pi/512
  assign cos2[6]  =  6'b001111;     //6pi/512
  assign sin2[7]  =  6'b111111;     //7pi/512
  assign cos2[7]  =  6'b001111;     //7pi/512
  assign sin2[8]  =  6'b111111;     //8pi/512
  assign cos2[8]  =  6'b001111;     //8pi/512
  assign sin2[9]  =  6'b111111;     //9pi/512
  assign cos2[9]  =  6'b001111;     //9pi/512
  assign sin2[10]  =  6'b111111;     //10pi/512
  assign cos2[10]  =  6'b001111;     //10pi/512
  assign sin2[11]  =  6'b111111;     //11pi/512
  assign cos2[11]  =  6'b001111;     //11pi/512
  assign sin2[12]  =  6'b111111;     //12pi/512
  assign cos2[12]  =  6'b001111;     //12pi/512
  assign sin2[13]  =  6'b111111;     //13pi/512
  assign cos2[13]  =  6'b001111;     //13pi/512
  assign sin2[14]  =  6'b111111;     //14pi/512
  assign cos2[14]  =  6'b001111;     //14pi/512
  assign sin2[15]  =  6'b111111;     //15pi/512
  assign cos2[15]  =  6'b001111;     //15pi/512
  assign sin2[16]  =  6'b111111;     //16pi/512
  assign cos2[16]  =  6'b001111;     //16pi/512
  assign sin2[17]  =  6'b111111;     //17pi/512
  assign cos2[17]  =  6'b001111;     //17pi/512
  assign sin2[18]  =  6'b111111;     //18pi/512
  assign cos2[18]  =  6'b001111;     //18pi/512
  assign sin2[19]  =  6'b111111;     //19pi/512
  assign cos2[19]  =  6'b001111;     //19pi/512
  assign sin2[20]  =  6'b111110;     //20pi/512
  assign cos2[20]  =  6'b001111;     //20pi/512
  assign sin2[21]  =  6'b111110;     //21pi/512
  assign cos2[21]  =  6'b001111;     //21pi/512
  assign sin2[22]  =  6'b111110;     //22pi/512
  assign cos2[22]  =  6'b001111;     //22pi/512
  assign sin2[23]  =  6'b111110;     //23pi/512
  assign cos2[23]  =  6'b001111;     //23pi/512
  assign sin2[24]  =  6'b111110;     //24pi/512
  assign cos2[24]  =  6'b001111;     //24pi/512
  assign sin2[25]  =  6'b111110;     //25pi/512
  assign cos2[25]  =  6'b001111;     //25pi/512
  assign sin2[26]  =  6'b111110;     //26pi/512
  assign cos2[26]  =  6'b001111;     //26pi/512
  assign sin2[27]  =  6'b111110;     //27pi/512
  assign cos2[27]  =  6'b001111;     //27pi/512
  assign sin2[28]  =  6'b111110;     //28pi/512
  assign cos2[28]  =  6'b001111;     //28pi/512
  assign sin2[29]  =  6'b111110;     //29pi/512
  assign cos2[29]  =  6'b001111;     //29pi/512
  assign sin2[30]  =  6'b111110;     //30pi/512
  assign cos2[30]  =  6'b001111;     //30pi/512
  assign sin2[31]  =  6'b111110;     //31pi/512
  assign cos2[31]  =  6'b001111;     //31pi/512
  assign sin2[32]  =  6'b111101;     //32pi/512
  assign cos2[32]  =  6'b001111;     //32pi/512
  assign sin2[33]  =  6'b111101;     //33pi/512
  assign cos2[33]  =  6'b001111;     //33pi/512
  assign sin2[34]  =  6'b111101;     //34pi/512
  assign cos2[34]  =  6'b001111;     //34pi/512
  assign sin2[35]  =  6'b111101;     //35pi/512
  assign cos2[35]  =  6'b001111;     //35pi/512
  assign sin2[36]  =  6'b111101;     //36pi/512
  assign cos2[36]  =  6'b001111;     //36pi/512
  assign sin2[37]  =  6'b111101;     //37pi/512
  assign cos2[37]  =  6'b001111;     //37pi/512
  assign sin2[38]  =  6'b111101;     //38pi/512
  assign cos2[38]  =  6'b001111;     //38pi/512
  assign sin2[39]  =  6'b111101;     //39pi/512
  assign cos2[39]  =  6'b001111;     //39pi/512
  assign sin2[40]  =  6'b111101;     //40pi/512
  assign cos2[40]  =  6'b001111;     //40pi/512
  assign sin2[41]  =  6'b111101;     //41pi/512
  assign cos2[41]  =  6'b001111;     //41pi/512
  assign sin2[42]  =  6'b111101;     //42pi/512
  assign cos2[42]  =  6'b001111;     //42pi/512
  assign sin2[43]  =  6'b111101;     //43pi/512
  assign cos2[43]  =  6'b001111;     //43pi/512
  assign sin2[44]  =  6'b111101;     //44pi/512
  assign cos2[44]  =  6'b001111;     //44pi/512
  assign sin2[45]  =  6'b111100;     //45pi/512
  assign cos2[45]  =  6'b001111;     //45pi/512
  assign sin2[46]  =  6'b111100;     //46pi/512
  assign cos2[46]  =  6'b001111;     //46pi/512
  assign sin2[47]  =  6'b111100;     //47pi/512
  assign cos2[47]  =  6'b001111;     //47pi/512
  assign sin2[48]  =  6'b111100;     //48pi/512
  assign cos2[48]  =  6'b001111;     //48pi/512
  assign sin2[49]  =  6'b111100;     //49pi/512
  assign cos2[49]  =  6'b001111;     //49pi/512
  assign sin2[50]  =  6'b111100;     //50pi/512
  assign cos2[50]  =  6'b001111;     //50pi/512
  assign sin2[51]  =  6'b111100;     //51pi/512
  assign cos2[51]  =  6'b001111;     //51pi/512
  assign sin2[52]  =  6'b111100;     //52pi/512
  assign cos2[52]  =  6'b001111;     //52pi/512
  assign sin2[53]  =  6'b111100;     //53pi/512
  assign cos2[53]  =  6'b001111;     //53pi/512
  assign sin2[54]  =  6'b111100;     //54pi/512
  assign cos2[54]  =  6'b001111;     //54pi/512
  assign sin2[55]  =  6'b111100;     //55pi/512
  assign cos2[55]  =  6'b001111;     //55pi/512
  assign sin2[56]  =  6'b111100;     //56pi/512
  assign cos2[56]  =  6'b001111;     //56pi/512
  assign sin2[57]  =  6'b111100;     //57pi/512
  assign cos2[57]  =  6'b001111;     //57pi/512
  assign sin2[58]  =  6'b111100;     //58pi/512
  assign cos2[58]  =  6'b001111;     //58pi/512
  assign sin2[59]  =  6'b111011;     //59pi/512
  assign cos2[59]  =  6'b001111;     //59pi/512
  assign sin2[60]  =  6'b111011;     //60pi/512
  assign cos2[60]  =  6'b001111;     //60pi/512
  assign sin2[61]  =  6'b111011;     //61pi/512
  assign cos2[61]  =  6'b001111;     //61pi/512
  assign sin2[62]  =  6'b111011;     //62pi/512
  assign cos2[62]  =  6'b001111;     //62pi/512
  assign sin2[63]  =  6'b111011;     //63pi/512
  assign cos2[63]  =  6'b001111;     //63pi/512
  assign sin2[64]  =  6'b111011;     //64pi/512
  assign cos2[64]  =  6'b001111;     //64pi/512
  assign sin2[65]  =  6'b111011;     //65pi/512
  assign cos2[65]  =  6'b001111;     //65pi/512
  assign sin2[66]  =  6'b111011;     //66pi/512
  assign cos2[66]  =  6'b001111;     //66pi/512
  assign sin2[67]  =  6'b111011;     //67pi/512
  assign cos2[67]  =  6'b001111;     //67pi/512
  assign sin2[68]  =  6'b111011;     //68pi/512
  assign cos2[68]  =  6'b001111;     //68pi/512
  assign sin2[69]  =  6'b111011;     //69pi/512
  assign cos2[69]  =  6'b001111;     //69pi/512
  assign sin2[70]  =  6'b111011;     //70pi/512
  assign cos2[70]  =  6'b001111;     //70pi/512
  assign sin2[71]  =  6'b111011;     //71pi/512
  assign cos2[71]  =  6'b001111;     //71pi/512
  assign sin2[72]  =  6'b111010;     //72pi/512
  assign cos2[72]  =  6'b001111;     //72pi/512
  assign sin2[73]  =  6'b111010;     //73pi/512
  assign cos2[73]  =  6'b001110;     //73pi/512
  assign sin2[74]  =  6'b111010;     //74pi/512
  assign cos2[74]  =  6'b001110;     //74pi/512
  assign sin2[75]  =  6'b111010;     //75pi/512
  assign cos2[75]  =  6'b001110;     //75pi/512
  assign sin2[76]  =  6'b111010;     //76pi/512
  assign cos2[76]  =  6'b001110;     //76pi/512
  assign sin2[77]  =  6'b111010;     //77pi/512
  assign cos2[77]  =  6'b001110;     //77pi/512
  assign sin2[78]  =  6'b111010;     //78pi/512
  assign cos2[78]  =  6'b001110;     //78pi/512
  assign sin2[79]  =  6'b111010;     //79pi/512
  assign cos2[79]  =  6'b001110;     //79pi/512
  assign sin2[80]  =  6'b111010;     //80pi/512
  assign cos2[80]  =  6'b001110;     //80pi/512
  assign sin2[81]  =  6'b111010;     //81pi/512
  assign cos2[81]  =  6'b001110;     //81pi/512
  assign sin2[82]  =  6'b111010;     //82pi/512
  assign cos2[82]  =  6'b001110;     //82pi/512
  assign sin2[83]  =  6'b111010;     //83pi/512
  assign cos2[83]  =  6'b001110;     //83pi/512
  assign sin2[84]  =  6'b111010;     //84pi/512
  assign cos2[84]  =  6'b001110;     //84pi/512
  assign sin2[85]  =  6'b111010;     //85pi/512
  assign cos2[85]  =  6'b001110;     //85pi/512
  assign sin2[86]  =  6'b111001;     //86pi/512
  assign cos2[86]  =  6'b001110;     //86pi/512
  assign sin2[87]  =  6'b111001;     //87pi/512
  assign cos2[87]  =  6'b001110;     //87pi/512
  assign sin2[88]  =  6'b111001;     //88pi/512
  assign cos2[88]  =  6'b001110;     //88pi/512
  assign sin2[89]  =  6'b111001;     //89pi/512
  assign cos2[89]  =  6'b001110;     //89pi/512
  assign sin2[90]  =  6'b111001;     //90pi/512
  assign cos2[90]  =  6'b001110;     //90pi/512
  assign sin2[91]  =  6'b111001;     //91pi/512
  assign cos2[91]  =  6'b001110;     //91pi/512
  assign sin2[92]  =  6'b111001;     //92pi/512
  assign cos2[92]  =  6'b001110;     //92pi/512
  assign sin2[93]  =  6'b111001;     //93pi/512
  assign cos2[93]  =  6'b001110;     //93pi/512
  assign sin2[94]  =  6'b111001;     //94pi/512
  assign cos2[94]  =  6'b001110;     //94pi/512
  assign sin2[95]  =  6'b111001;     //95pi/512
  assign cos2[95]  =  6'b001110;     //95pi/512
  assign sin2[96]  =  6'b111001;     //96pi/512
  assign cos2[96]  =  6'b001110;     //96pi/512
  assign sin2[97]  =  6'b111001;     //97pi/512
  assign cos2[97]  =  6'b001110;     //97pi/512
  assign sin2[98]  =  6'b111001;     //98pi/512
  assign cos2[98]  =  6'b001110;     //98pi/512
  assign sin2[99]  =  6'b111001;     //99pi/512
  assign cos2[99]  =  6'b001110;     //99pi/512
  assign sin2[100]  =  6'b111000;     //100pi/512
  assign cos2[100]  =  6'b001110;     //100pi/512
  assign sin2[101]  =  6'b111000;     //101pi/512
  assign cos2[101]  =  6'b001110;     //101pi/512
  assign sin2[102]  =  6'b111000;     //102pi/512
  assign cos2[102]  =  6'b001110;     //102pi/512
  assign sin2[103]  =  6'b111000;     //103pi/512
  assign cos2[103]  =  6'b001101;     //103pi/512
  assign sin2[104]  =  6'b111000;     //104pi/512
  assign cos2[104]  =  6'b001101;     //104pi/512
  assign sin2[105]  =  6'b111000;     //105pi/512
  assign cos2[105]  =  6'b001101;     //105pi/512
  assign sin2[106]  =  6'b111000;     //106pi/512
  assign cos2[106]  =  6'b001101;     //106pi/512
  assign sin2[107]  =  6'b111000;     //107pi/512
  assign cos2[107]  =  6'b001101;     //107pi/512
  assign sin2[108]  =  6'b111000;     //108pi/512
  assign cos2[108]  =  6'b001101;     //108pi/512
  assign sin2[109]  =  6'b111000;     //109pi/512
  assign cos2[109]  =  6'b001101;     //109pi/512
  assign sin2[110]  =  6'b111000;     //110pi/512
  assign cos2[110]  =  6'b001101;     //110pi/512
  assign sin2[111]  =  6'b111000;     //111pi/512
  assign cos2[111]  =  6'b001101;     //111pi/512
  assign sin2[112]  =  6'b111000;     //112pi/512
  assign cos2[112]  =  6'b001101;     //112pi/512
  assign sin2[113]  =  6'b111000;     //113pi/512
  assign cos2[113]  =  6'b001101;     //113pi/512
  assign sin2[114]  =  6'b111000;     //114pi/512
  assign cos2[114]  =  6'b001101;     //114pi/512
  assign sin2[115]  =  6'b110111;     //115pi/512
  assign cos2[115]  =  6'b001101;     //115pi/512
  assign sin2[116]  =  6'b110111;     //116pi/512
  assign cos2[116]  =  6'b001101;     //116pi/512
  assign sin2[117]  =  6'b110111;     //117pi/512
  assign cos2[117]  =  6'b001101;     //117pi/512
  assign sin2[118]  =  6'b110111;     //118pi/512
  assign cos2[118]  =  6'b001101;     //118pi/512
  assign sin2[119]  =  6'b110111;     //119pi/512
  assign cos2[119]  =  6'b001101;     //119pi/512
  assign sin2[120]  =  6'b110111;     //120pi/512
  assign cos2[120]  =  6'b001101;     //120pi/512
  assign sin2[121]  =  6'b110111;     //121pi/512
  assign cos2[121]  =  6'b001101;     //121pi/512
  assign sin2[122]  =  6'b110111;     //122pi/512
  assign cos2[122]  =  6'b001101;     //122pi/512
  assign sin2[123]  =  6'b110111;     //123pi/512
  assign cos2[123]  =  6'b001101;     //123pi/512
  assign sin2[124]  =  6'b110111;     //124pi/512
  assign cos2[124]  =  6'b001101;     //124pi/512
  assign sin2[125]  =  6'b110111;     //125pi/512
  assign cos2[125]  =  6'b001101;     //125pi/512
  assign sin2[126]  =  6'b110111;     //126pi/512
  assign cos2[126]  =  6'b001101;     //126pi/512
  assign sin2[127]  =  6'b110111;     //127pi/512
  assign cos2[127]  =  6'b001100;     //127pi/512
  assign sin2[128]  =  6'b110111;     //128pi/512
  assign cos2[128]  =  6'b001100;     //128pi/512
  assign sin2[129]  =  6'b110111;     //129pi/512
  assign cos2[129]  =  6'b001100;     //129pi/512
  assign sin2[130]  =  6'b110110;     //130pi/512
  assign cos2[130]  =  6'b001100;     //130pi/512
  assign sin2[131]  =  6'b110110;     //131pi/512
  assign cos2[131]  =  6'b001100;     //131pi/512
  assign sin2[132]  =  6'b110110;     //132pi/512
  assign cos2[132]  =  6'b001100;     //132pi/512
  assign sin2[133]  =  6'b110110;     //133pi/512
  assign cos2[133]  =  6'b001100;     //133pi/512
  assign sin2[134]  =  6'b110110;     //134pi/512
  assign cos2[134]  =  6'b001100;     //134pi/512
  assign sin2[135]  =  6'b110110;     //135pi/512
  assign cos2[135]  =  6'b001100;     //135pi/512
  assign sin2[136]  =  6'b110110;     //136pi/512
  assign cos2[136]  =  6'b001100;     //136pi/512
  assign sin2[137]  =  6'b110110;     //137pi/512
  assign cos2[137]  =  6'b001100;     //137pi/512
  assign sin2[138]  =  6'b110110;     //138pi/512
  assign cos2[138]  =  6'b001100;     //138pi/512
  assign sin2[139]  =  6'b110110;     //139pi/512
  assign cos2[139]  =  6'b001100;     //139pi/512
  assign sin2[140]  =  6'b110110;     //140pi/512
  assign cos2[140]  =  6'b001100;     //140pi/512
  assign sin2[141]  =  6'b110110;     //141pi/512
  assign cos2[141]  =  6'b001100;     //141pi/512
  assign sin2[142]  =  6'b110110;     //142pi/512
  assign cos2[142]  =  6'b001100;     //142pi/512
  assign sin2[143]  =  6'b110110;     //143pi/512
  assign cos2[143]  =  6'b001100;     //143pi/512
  assign sin2[144]  =  6'b110110;     //144pi/512
  assign cos2[144]  =  6'b001100;     //144pi/512
  assign sin2[145]  =  6'b110110;     //145pi/512
  assign cos2[145]  =  6'b001100;     //145pi/512
  assign sin2[146]  =  6'b110101;     //146pi/512
  assign cos2[146]  =  6'b001100;     //146pi/512
  assign sin2[147]  =  6'b110101;     //147pi/512
  assign cos2[147]  =  6'b001100;     //147pi/512
  assign sin2[148]  =  6'b110101;     //148pi/512
  assign cos2[148]  =  6'b001011;     //148pi/512
  assign sin2[149]  =  6'b110101;     //149pi/512
  assign cos2[149]  =  6'b001011;     //149pi/512
  assign sin2[150]  =  6'b110101;     //150pi/512
  assign cos2[150]  =  6'b001011;     //150pi/512
  assign sin2[151]  =  6'b110101;     //151pi/512
  assign cos2[151]  =  6'b001011;     //151pi/512
  assign sin2[152]  =  6'b110101;     //152pi/512
  assign cos2[152]  =  6'b001011;     //152pi/512
  assign sin2[153]  =  6'b110101;     //153pi/512
  assign cos2[153]  =  6'b001011;     //153pi/512
  assign sin2[154]  =  6'b110101;     //154pi/512
  assign cos2[154]  =  6'b001011;     //154pi/512
  assign sin2[155]  =  6'b110101;     //155pi/512
  assign cos2[155]  =  6'b001011;     //155pi/512
  assign sin2[156]  =  6'b110101;     //156pi/512
  assign cos2[156]  =  6'b001011;     //156pi/512
  assign sin2[157]  =  6'b110101;     //157pi/512
  assign cos2[157]  =  6'b001011;     //157pi/512
  assign sin2[158]  =  6'b110101;     //158pi/512
  assign cos2[158]  =  6'b001011;     //158pi/512
  assign sin2[159]  =  6'b110101;     //159pi/512
  assign cos2[159]  =  6'b001011;     //159pi/512
  assign sin2[160]  =  6'b110101;     //160pi/512
  assign cos2[160]  =  6'b001011;     //160pi/512
  assign sin2[161]  =  6'b110101;     //161pi/512
  assign cos2[161]  =  6'b001011;     //161pi/512
  assign sin2[162]  =  6'b110101;     //162pi/512
  assign cos2[162]  =  6'b001011;     //162pi/512
  assign sin2[163]  =  6'b110101;     //163pi/512
  assign cos2[163]  =  6'b001011;     //163pi/512
  assign sin2[164]  =  6'b110100;     //164pi/512
  assign cos2[164]  =  6'b001011;     //164pi/512
  assign sin2[165]  =  6'b110100;     //165pi/512
  assign cos2[165]  =  6'b001011;     //165pi/512
  assign sin2[166]  =  6'b110100;     //166pi/512
  assign cos2[166]  =  6'b001010;     //166pi/512
  assign sin2[167]  =  6'b110100;     //167pi/512
  assign cos2[167]  =  6'b001010;     //167pi/512
  assign sin2[168]  =  6'b110100;     //168pi/512
  assign cos2[168]  =  6'b001010;     //168pi/512
  assign sin2[169]  =  6'b110100;     //169pi/512
  assign cos2[169]  =  6'b001010;     //169pi/512
  assign sin2[170]  =  6'b110100;     //170pi/512
  assign cos2[170]  =  6'b001010;     //170pi/512
  assign sin2[171]  =  6'b110100;     //171pi/512
  assign cos2[171]  =  6'b001010;     //171pi/512
  assign sin2[172]  =  6'b110100;     //172pi/512
  assign cos2[172]  =  6'b001010;     //172pi/512
  assign sin2[173]  =  6'b110100;     //173pi/512
  assign cos2[173]  =  6'b001010;     //173pi/512
  assign sin2[174]  =  6'b110100;     //174pi/512
  assign cos2[174]  =  6'b001010;     //174pi/512
  assign sin2[175]  =  6'b110100;     //175pi/512
  assign cos2[175]  =  6'b001010;     //175pi/512
  assign sin2[176]  =  6'b110100;     //176pi/512
  assign cos2[176]  =  6'b001010;     //176pi/512
  assign sin2[177]  =  6'b110100;     //177pi/512
  assign cos2[177]  =  6'b001010;     //177pi/512
  assign sin2[178]  =  6'b110100;     //178pi/512
  assign cos2[178]  =  6'b001010;     //178pi/512
  assign sin2[179]  =  6'b110100;     //179pi/512
  assign cos2[179]  =  6'b001010;     //179pi/512
  assign sin2[180]  =  6'b110100;     //180pi/512
  assign cos2[180]  =  6'b001010;     //180pi/512
  assign sin2[181]  =  6'b110100;     //181pi/512
  assign cos2[181]  =  6'b001010;     //181pi/512
  assign sin2[182]  =  6'b110100;     //182pi/512
  assign cos2[182]  =  6'b001010;     //182pi/512
  assign sin2[183]  =  6'b110011;     //183pi/512
  assign cos2[183]  =  6'b001001;     //183pi/512
  assign sin2[184]  =  6'b110011;     //184pi/512
  assign cos2[184]  =  6'b001001;     //184pi/512
  assign sin2[185]  =  6'b110011;     //185pi/512
  assign cos2[185]  =  6'b001001;     //185pi/512
  assign sin2[186]  =  6'b110011;     //186pi/512
  assign cos2[186]  =  6'b001001;     //186pi/512
  assign sin2[187]  =  6'b110011;     //187pi/512
  assign cos2[187]  =  6'b001001;     //187pi/512
  assign sin2[188]  =  6'b110011;     //188pi/512
  assign cos2[188]  =  6'b001001;     //188pi/512
  assign sin2[189]  =  6'b110011;     //189pi/512
  assign cos2[189]  =  6'b001001;     //189pi/512
  assign sin2[190]  =  6'b110011;     //190pi/512
  assign cos2[190]  =  6'b001001;     //190pi/512
  assign sin2[191]  =  6'b110011;     //191pi/512
  assign cos2[191]  =  6'b001001;     //191pi/512
  assign sin2[192]  =  6'b110011;     //192pi/512
  assign cos2[192]  =  6'b001001;     //192pi/512
  assign sin2[193]  =  6'b110011;     //193pi/512
  assign cos2[193]  =  6'b001001;     //193pi/512
  assign sin2[194]  =  6'b110011;     //194pi/512
  assign cos2[194]  =  6'b001001;     //194pi/512
  assign sin2[195]  =  6'b110011;     //195pi/512
  assign cos2[195]  =  6'b001001;     //195pi/512
  assign sin2[196]  =  6'b110011;     //196pi/512
  assign cos2[196]  =  6'b001001;     //196pi/512
  assign sin2[197]  =  6'b110011;     //197pi/512
  assign cos2[197]  =  6'b001001;     //197pi/512
  assign sin2[198]  =  6'b110011;     //198pi/512
  assign cos2[198]  =  6'b001001;     //198pi/512
  assign sin2[199]  =  6'b110011;     //199pi/512
  assign cos2[199]  =  6'b001000;     //199pi/512
  assign sin2[200]  =  6'b110011;     //200pi/512
  assign cos2[200]  =  6'b001000;     //200pi/512
  assign sin2[201]  =  6'b110011;     //201pi/512
  assign cos2[201]  =  6'b001000;     //201pi/512
  assign sin2[202]  =  6'b110011;     //202pi/512
  assign cos2[202]  =  6'b001000;     //202pi/512
  assign sin2[203]  =  6'b110011;     //203pi/512
  assign cos2[203]  =  6'b001000;     //203pi/512
  assign sin2[204]  =  6'b110011;     //204pi/512
  assign cos2[204]  =  6'b001000;     //204pi/512
  assign sin2[205]  =  6'b110010;     //205pi/512
  assign cos2[205]  =  6'b001000;     //205pi/512
  assign sin2[206]  =  6'b110010;     //206pi/512
  assign cos2[206]  =  6'b001000;     //206pi/512
  assign sin2[207]  =  6'b110010;     //207pi/512
  assign cos2[207]  =  6'b001000;     //207pi/512
  assign sin2[208]  =  6'b110010;     //208pi/512
  assign cos2[208]  =  6'b001000;     //208pi/512
  assign sin2[209]  =  6'b110010;     //209pi/512
  assign cos2[209]  =  6'b001000;     //209pi/512
  assign sin2[210]  =  6'b110010;     //210pi/512
  assign cos2[210]  =  6'b001000;     //210pi/512
  assign sin2[211]  =  6'b110010;     //211pi/512
  assign cos2[211]  =  6'b001000;     //211pi/512
  assign sin2[212]  =  6'b110010;     //212pi/512
  assign cos2[212]  =  6'b001000;     //212pi/512
  assign sin2[213]  =  6'b110010;     //213pi/512
  assign cos2[213]  =  6'b001000;     //213pi/512
  assign sin2[214]  =  6'b110010;     //214pi/512
  assign cos2[214]  =  6'b000111;     //214pi/512
  assign sin2[215]  =  6'b110010;     //215pi/512
  assign cos2[215]  =  6'b000111;     //215pi/512
  assign sin2[216]  =  6'b110010;     //216pi/512
  assign cos2[216]  =  6'b000111;     //216pi/512
  assign sin2[217]  =  6'b110010;     //217pi/512
  assign cos2[217]  =  6'b000111;     //217pi/512
  assign sin2[218]  =  6'b110010;     //218pi/512
  assign cos2[218]  =  6'b000111;     //218pi/512
  assign sin2[219]  =  6'b110010;     //219pi/512
  assign cos2[219]  =  6'b000111;     //219pi/512
  assign sin2[220]  =  6'b110010;     //220pi/512
  assign cos2[220]  =  6'b000111;     //220pi/512
  assign sin2[221]  =  6'b110010;     //221pi/512
  assign cos2[221]  =  6'b000111;     //221pi/512
  assign sin2[222]  =  6'b110010;     //222pi/512
  assign cos2[222]  =  6'b000111;     //222pi/512
  assign sin2[223]  =  6'b110010;     //223pi/512
  assign cos2[223]  =  6'b000111;     //223pi/512
  assign sin2[224]  =  6'b110010;     //224pi/512
  assign cos2[224]  =  6'b000111;     //224pi/512
  assign sin2[225]  =  6'b110010;     //225pi/512
  assign cos2[225]  =  6'b000111;     //225pi/512
  assign sin2[226]  =  6'b110010;     //226pi/512
  assign cos2[226]  =  6'b000111;     //226pi/512
  assign sin2[227]  =  6'b110010;     //227pi/512
  assign cos2[227]  =  6'b000111;     //227pi/512
  assign sin2[228]  =  6'b110010;     //228pi/512
  assign cos2[228]  =  6'b000110;     //228pi/512
  assign sin2[229]  =  6'b110010;     //229pi/512
  assign cos2[229]  =  6'b000110;     //229pi/512
  assign sin2[230]  =  6'b110010;     //230pi/512
  assign cos2[230]  =  6'b000110;     //230pi/512
  assign sin2[231]  =  6'b110010;     //231pi/512
  assign cos2[231]  =  6'b000110;     //231pi/512
  assign sin2[232]  =  6'b110001;     //232pi/512
  assign cos2[232]  =  6'b000110;     //232pi/512
  assign sin2[233]  =  6'b110001;     //233pi/512
  assign cos2[233]  =  6'b000110;     //233pi/512
  assign sin2[234]  =  6'b110001;     //234pi/512
  assign cos2[234]  =  6'b000110;     //234pi/512
  assign sin2[235]  =  6'b110001;     //235pi/512
  assign cos2[235]  =  6'b000110;     //235pi/512
  assign sin2[236]  =  6'b110001;     //236pi/512
  assign cos2[236]  =  6'b000110;     //236pi/512
  assign sin2[237]  =  6'b110001;     //237pi/512
  assign cos2[237]  =  6'b000110;     //237pi/512
  assign sin2[238]  =  6'b110001;     //238pi/512
  assign cos2[238]  =  6'b000110;     //238pi/512
  assign sin2[239]  =  6'b110001;     //239pi/512
  assign cos2[239]  =  6'b000110;     //239pi/512
  assign sin2[240]  =  6'b110001;     //240pi/512
  assign cos2[240]  =  6'b000110;     //240pi/512
  assign sin2[241]  =  6'b110001;     //241pi/512
  assign cos2[241]  =  6'b000110;     //241pi/512
  assign sin2[242]  =  6'b110001;     //242pi/512
  assign cos2[242]  =  6'b000101;     //242pi/512
  assign sin2[243]  =  6'b110001;     //243pi/512
  assign cos2[243]  =  6'b000101;     //243pi/512
  assign sin2[244]  =  6'b110001;     //244pi/512
  assign cos2[244]  =  6'b000101;     //244pi/512
  assign sin2[245]  =  6'b110001;     //245pi/512
  assign cos2[245]  =  6'b000101;     //245pi/512
  assign sin2[246]  =  6'b110001;     //246pi/512
  assign cos2[246]  =  6'b000101;     //246pi/512
  assign sin2[247]  =  6'b110001;     //247pi/512
  assign cos2[247]  =  6'b000101;     //247pi/512
  assign sin2[248]  =  6'b110001;     //248pi/512
  assign cos2[248]  =  6'b000101;     //248pi/512
  assign sin2[249]  =  6'b110001;     //249pi/512
  assign cos2[249]  =  6'b000101;     //249pi/512
  assign sin2[250]  =  6'b110001;     //250pi/512
  assign cos2[250]  =  6'b000101;     //250pi/512
  assign sin2[251]  =  6'b110001;     //251pi/512
  assign cos2[251]  =  6'b000101;     //251pi/512
  assign sin2[252]  =  6'b110001;     //252pi/512
  assign cos2[252]  =  6'b000101;     //252pi/512
  assign sin2[253]  =  6'b110001;     //253pi/512
  assign cos2[253]  =  6'b000101;     //253pi/512
  assign sin2[254]  =  6'b110001;     //254pi/512
  assign cos2[254]  =  6'b000101;     //254pi/512
  assign sin2[255]  =  6'b110001;     //255pi/512
  assign cos2[255]  =  6'b000101;     //255pi/512
  assign sin2[256]  =  6'b110001;     //256pi/512
  assign cos2[256]  =  6'b000100;     //256pi/512
  assign sin2[257]  =  6'b110001;     //257pi/512
  assign cos2[257]  =  6'b000100;     //257pi/512
  assign sin2[258]  =  6'b110001;     //258pi/512
  assign cos2[258]  =  6'b000100;     //258pi/512
  assign sin2[259]  =  6'b110001;     //259pi/512
  assign cos2[259]  =  6'b000100;     //259pi/512
  assign sin2[260]  =  6'b110001;     //260pi/512
  assign cos2[260]  =  6'b000100;     //260pi/512
  assign sin2[261]  =  6'b110001;     //261pi/512
  assign cos2[261]  =  6'b000100;     //261pi/512
  assign sin2[262]  =  6'b110001;     //262pi/512
  assign cos2[262]  =  6'b000100;     //262pi/512
  assign sin2[263]  =  6'b110001;     //263pi/512
  assign cos2[263]  =  6'b000100;     //263pi/512
  assign sin2[264]  =  6'b110001;     //264pi/512
  assign cos2[264]  =  6'b000100;     //264pi/512
  assign sin2[265]  =  6'b110001;     //265pi/512
  assign cos2[265]  =  6'b000100;     //265pi/512
  assign sin2[266]  =  6'b110001;     //266pi/512
  assign cos2[266]  =  6'b000100;     //266pi/512
  assign sin2[267]  =  6'b110001;     //267pi/512
  assign cos2[267]  =  6'b000100;     //267pi/512
  assign sin2[268]  =  6'b110001;     //268pi/512
  assign cos2[268]  =  6'b000100;     //268pi/512
  assign sin2[269]  =  6'b110000;     //269pi/512
  assign cos2[269]  =  6'b000011;     //269pi/512
  assign sin2[270]  =  6'b110000;     //270pi/512
  assign cos2[270]  =  6'b000011;     //270pi/512
  assign sin2[271]  =  6'b110000;     //271pi/512
  assign cos2[271]  =  6'b000011;     //271pi/512
  assign sin2[272]  =  6'b110000;     //272pi/512
  assign cos2[272]  =  6'b000011;     //272pi/512
  assign sin2[273]  =  6'b110000;     //273pi/512
  assign cos2[273]  =  6'b000011;     //273pi/512
  assign sin2[274]  =  6'b110000;     //274pi/512
  assign cos2[274]  =  6'b000011;     //274pi/512
  assign sin2[275]  =  6'b110000;     //275pi/512
  assign cos2[275]  =  6'b000011;     //275pi/512
  assign sin2[276]  =  6'b110000;     //276pi/512
  assign cos2[276]  =  6'b000011;     //276pi/512
  assign sin2[277]  =  6'b110000;     //277pi/512
  assign cos2[277]  =  6'b000011;     //277pi/512
  assign sin2[278]  =  6'b110000;     //278pi/512
  assign cos2[278]  =  6'b000011;     //278pi/512
  assign sin2[279]  =  6'b110000;     //279pi/512
  assign cos2[279]  =  6'b000011;     //279pi/512
  assign sin2[280]  =  6'b110000;     //280pi/512
  assign cos2[280]  =  6'b000011;     //280pi/512
  assign sin2[281]  =  6'b110000;     //281pi/512
  assign cos2[281]  =  6'b000011;     //281pi/512
  assign sin2[282]  =  6'b110000;     //282pi/512
  assign cos2[282]  =  6'b000010;     //282pi/512
  assign sin2[283]  =  6'b110000;     //283pi/512
  assign cos2[283]  =  6'b000010;     //283pi/512
  assign sin2[284]  =  6'b110000;     //284pi/512
  assign cos2[284]  =  6'b000010;     //284pi/512
  assign sin2[285]  =  6'b110000;     //285pi/512
  assign cos2[285]  =  6'b000010;     //285pi/512
  assign sin2[286]  =  6'b110000;     //286pi/512
  assign cos2[286]  =  6'b000010;     //286pi/512
  assign sin2[287]  =  6'b110000;     //287pi/512
  assign cos2[287]  =  6'b000010;     //287pi/512
  assign sin2[288]  =  6'b110000;     //288pi/512
  assign cos2[288]  =  6'b000010;     //288pi/512
  assign sin2[289]  =  6'b110000;     //289pi/512
  assign cos2[289]  =  6'b000010;     //289pi/512
  assign sin2[290]  =  6'b110000;     //290pi/512
  assign cos2[290]  =  6'b000010;     //290pi/512
  assign sin2[291]  =  6'b110000;     //291pi/512
  assign cos2[291]  =  6'b000010;     //291pi/512
  assign sin2[292]  =  6'b110000;     //292pi/512
  assign cos2[292]  =  6'b000010;     //292pi/512
  assign sin2[293]  =  6'b110000;     //293pi/512
  assign cos2[293]  =  6'b000010;     //293pi/512
  assign sin2[294]  =  6'b110000;     //294pi/512
  assign cos2[294]  =  6'b000010;     //294pi/512
  assign sin2[295]  =  6'b110000;     //295pi/512
  assign cos2[295]  =  6'b000001;     //295pi/512
  assign sin2[296]  =  6'b110000;     //296pi/512
  assign cos2[296]  =  6'b000001;     //296pi/512
  assign sin2[297]  =  6'b110000;     //297pi/512
  assign cos2[297]  =  6'b000001;     //297pi/512
  assign sin2[298]  =  6'b110000;     //298pi/512
  assign cos2[298]  =  6'b000001;     //298pi/512
  assign sin2[299]  =  6'b110000;     //299pi/512
  assign cos2[299]  =  6'b000001;     //299pi/512
  assign sin2[300]  =  6'b110000;     //300pi/512
  assign cos2[300]  =  6'b000001;     //300pi/512
  assign sin2[301]  =  6'b110000;     //301pi/512
  assign cos2[301]  =  6'b000001;     //301pi/512
  assign sin2[302]  =  6'b110000;     //302pi/512
  assign cos2[302]  =  6'b000001;     //302pi/512
  assign sin2[303]  =  6'b110000;     //303pi/512
  assign cos2[303]  =  6'b000001;     //303pi/512
  assign sin2[304]  =  6'b110000;     //304pi/512
  assign cos2[304]  =  6'b000001;     //304pi/512
  assign sin2[305]  =  6'b110000;     //305pi/512
  assign cos2[305]  =  6'b000001;     //305pi/512
  assign sin2[306]  =  6'b110000;     //306pi/512
  assign cos2[306]  =  6'b000001;     //306pi/512
  assign sin2[307]  =  6'b110000;     //307pi/512
  assign cos2[307]  =  6'b000001;     //307pi/512
  assign sin2[308]  =  6'b110000;     //308pi/512
  assign cos2[308]  =  6'b000000;     //308pi/512
  assign sin2[309]  =  6'b110000;     //309pi/512
  assign cos2[309]  =  6'b000000;     //309pi/512
  assign sin2[310]  =  6'b110000;     //310pi/512
  assign cos2[310]  =  6'b000000;     //310pi/512
  assign sin2[311]  =  6'b110000;     //311pi/512
  assign cos2[311]  =  6'b000000;     //311pi/512
  assign sin2[312]  =  6'b110000;     //312pi/512
  assign cos2[312]  =  6'b000000;     //312pi/512
  assign sin2[313]  =  6'b110000;     //313pi/512
  assign cos2[313]  =  6'b000000;     //313pi/512
  assign sin2[314]  =  6'b110000;     //314pi/512
  assign cos2[314]  =  6'b000000;     //314pi/512
  assign sin2[315]  =  6'b110000;     //315pi/512
  assign cos2[315]  =  6'b000000;     //315pi/512
  assign sin2[316]  =  6'b110000;     //316pi/512
  assign cos2[316]  =  6'b000000;     //316pi/512
  assign sin2[317]  =  6'b110000;     //317pi/512
  assign cos2[317]  =  6'b000000;     //317pi/512
  assign sin2[318]  =  6'b110000;     //318pi/512
  assign cos2[318]  =  6'b000000;     //318pi/512
  assign sin2[319]  =  6'b110000;     //319pi/512
  assign cos2[319]  =  6'b000000;     //319pi/512
  assign sin2[320]  =  6'b110000;     //320pi/512
  assign cos2[320]  =  6'b000000;     //320pi/512
  assign sin2[321]  =  6'b110000;     //321pi/512
  assign cos2[321]  =  6'b000000;     //321pi/512
  assign sin2[322]  =  6'b110000;     //322pi/512
  assign cos2[322]  =  6'b000000;     //322pi/512
  assign sin2[323]  =  6'b110000;     //323pi/512
  assign cos2[323]  =  6'b000000;     //323pi/512
  assign sin2[324]  =  6'b110000;     //324pi/512
  assign cos2[324]  =  6'b000000;     //324pi/512
  assign sin2[325]  =  6'b110000;     //325pi/512
  assign cos2[325]  =  6'b000000;     //325pi/512
  assign sin2[326]  =  6'b110000;     //326pi/512
  assign cos2[326]  =  6'b000000;     //326pi/512
  assign sin2[327]  =  6'b110000;     //327pi/512
  assign cos2[327]  =  6'b111111;     //327pi/512
  assign sin2[328]  =  6'b110000;     //328pi/512
  assign cos2[328]  =  6'b111111;     //328pi/512
  assign sin2[329]  =  6'b110000;     //329pi/512
  assign cos2[329]  =  6'b111111;     //329pi/512
  assign sin2[330]  =  6'b110000;     //330pi/512
  assign cos2[330]  =  6'b111111;     //330pi/512
  assign sin2[331]  =  6'b110000;     //331pi/512
  assign cos2[331]  =  6'b111111;     //331pi/512
  assign sin2[332]  =  6'b110000;     //332pi/512
  assign cos2[332]  =  6'b111111;     //332pi/512
  assign sin2[333]  =  6'b110000;     //333pi/512
  assign cos2[333]  =  6'b111111;     //333pi/512
  assign sin2[334]  =  6'b110000;     //334pi/512
  assign cos2[334]  =  6'b111111;     //334pi/512
  assign sin2[335]  =  6'b110000;     //335pi/512
  assign cos2[335]  =  6'b111111;     //335pi/512
  assign sin2[336]  =  6'b110000;     //336pi/512
  assign cos2[336]  =  6'b111111;     //336pi/512
  assign sin2[337]  =  6'b110000;     //337pi/512
  assign cos2[337]  =  6'b111111;     //337pi/512
  assign sin2[338]  =  6'b110000;     //338pi/512
  assign cos2[338]  =  6'b111111;     //338pi/512
  assign sin2[339]  =  6'b110000;     //339pi/512
  assign cos2[339]  =  6'b111111;     //339pi/512
  assign sin2[340]  =  6'b110000;     //340pi/512
  assign cos2[340]  =  6'b111110;     //340pi/512
  assign sin2[341]  =  6'b110000;     //341pi/512
  assign cos2[341]  =  6'b111110;     //341pi/512
  assign sin2[342]  =  6'b110000;     //342pi/512
  assign cos2[342]  =  6'b111110;     //342pi/512
  assign sin2[343]  =  6'b110000;     //343pi/512
  assign cos2[343]  =  6'b111110;     //343pi/512
  assign sin2[344]  =  6'b110000;     //344pi/512
  assign cos2[344]  =  6'b111110;     //344pi/512
  assign sin2[345]  =  6'b110000;     //345pi/512
  assign cos2[345]  =  6'b111110;     //345pi/512
  assign sin2[346]  =  6'b110000;     //346pi/512
  assign cos2[346]  =  6'b111110;     //346pi/512
  assign sin2[347]  =  6'b110000;     //347pi/512
  assign cos2[347]  =  6'b111110;     //347pi/512
  assign sin2[348]  =  6'b110000;     //348pi/512
  assign cos2[348]  =  6'b111110;     //348pi/512
  assign sin2[349]  =  6'b110000;     //349pi/512
  assign cos2[349]  =  6'b111110;     //349pi/512
  assign sin2[350]  =  6'b110000;     //350pi/512
  assign cos2[350]  =  6'b111110;     //350pi/512
  assign sin2[351]  =  6'b110000;     //351pi/512
  assign cos2[351]  =  6'b111110;     //351pi/512
  assign sin2[352]  =  6'b110000;     //352pi/512
  assign cos2[352]  =  6'b111101;     //352pi/512
  assign sin2[353]  =  6'b110000;     //353pi/512
  assign cos2[353]  =  6'b111101;     //353pi/512
  assign sin2[354]  =  6'b110000;     //354pi/512
  assign cos2[354]  =  6'b111101;     //354pi/512
  assign sin2[355]  =  6'b110000;     //355pi/512
  assign cos2[355]  =  6'b111101;     //355pi/512
  assign sin2[356]  =  6'b110000;     //356pi/512
  assign cos2[356]  =  6'b111101;     //356pi/512
  assign sin2[357]  =  6'b110000;     //357pi/512
  assign cos2[357]  =  6'b111101;     //357pi/512
  assign sin2[358]  =  6'b110000;     //358pi/512
  assign cos2[358]  =  6'b111101;     //358pi/512
  assign sin2[359]  =  6'b110000;     //359pi/512
  assign cos2[359]  =  6'b111101;     //359pi/512
  assign sin2[360]  =  6'b110000;     //360pi/512
  assign cos2[360]  =  6'b111101;     //360pi/512
  assign sin2[361]  =  6'b110000;     //361pi/512
  assign cos2[361]  =  6'b111101;     //361pi/512
  assign sin2[362]  =  6'b110000;     //362pi/512
  assign cos2[362]  =  6'b111101;     //362pi/512
  assign sin2[363]  =  6'b110000;     //363pi/512
  assign cos2[363]  =  6'b111101;     //363pi/512
  assign sin2[364]  =  6'b110000;     //364pi/512
  assign cos2[364]  =  6'b111101;     //364pi/512
  assign sin2[365]  =  6'b110000;     //365pi/512
  assign cos2[365]  =  6'b111100;     //365pi/512
  assign sin2[366]  =  6'b110000;     //366pi/512
  assign cos2[366]  =  6'b111100;     //366pi/512
  assign sin2[367]  =  6'b110000;     //367pi/512
  assign cos2[367]  =  6'b111100;     //367pi/512
  assign sin2[368]  =  6'b110000;     //368pi/512
  assign cos2[368]  =  6'b111100;     //368pi/512
  assign sin2[369]  =  6'b110000;     //369pi/512
  assign cos2[369]  =  6'b111100;     //369pi/512
  assign sin2[370]  =  6'b110000;     //370pi/512
  assign cos2[370]  =  6'b111100;     //370pi/512
  assign sin2[371]  =  6'b110000;     //371pi/512
  assign cos2[371]  =  6'b111100;     //371pi/512
  assign sin2[372]  =  6'b110001;     //372pi/512
  assign cos2[372]  =  6'b111100;     //372pi/512
  assign sin2[373]  =  6'b110001;     //373pi/512
  assign cos2[373]  =  6'b111100;     //373pi/512
  assign sin2[374]  =  6'b110001;     //374pi/512
  assign cos2[374]  =  6'b111100;     //374pi/512
  assign sin2[375]  =  6'b110001;     //375pi/512
  assign cos2[375]  =  6'b111100;     //375pi/512
  assign sin2[376]  =  6'b110001;     //376pi/512
  assign cos2[376]  =  6'b111100;     //376pi/512
  assign sin2[377]  =  6'b110001;     //377pi/512
  assign cos2[377]  =  6'b111100;     //377pi/512
  assign sin2[378]  =  6'b110001;     //378pi/512
  assign cos2[378]  =  6'b111100;     //378pi/512
  assign sin2[379]  =  6'b110001;     //379pi/512
  assign cos2[379]  =  6'b111011;     //379pi/512
  assign sin2[380]  =  6'b110001;     //380pi/512
  assign cos2[380]  =  6'b111011;     //380pi/512
  assign sin2[381]  =  6'b110001;     //381pi/512
  assign cos2[381]  =  6'b111011;     //381pi/512
  assign sin2[382]  =  6'b110001;     //382pi/512
  assign cos2[382]  =  6'b111011;     //382pi/512
  assign sin2[383]  =  6'b110001;     //383pi/512
  assign cos2[383]  =  6'b111011;     //383pi/512
  assign sin2[384]  =  6'b110001;     //384pi/512
  assign cos2[384]  =  6'b111011;     //384pi/512
  assign sin2[385]  =  6'b110001;     //385pi/512
  assign cos2[385]  =  6'b111011;     //385pi/512
  assign sin2[386]  =  6'b110001;     //386pi/512
  assign cos2[386]  =  6'b111011;     //386pi/512
  assign sin2[387]  =  6'b110001;     //387pi/512
  assign cos2[387]  =  6'b111011;     //387pi/512
  assign sin2[388]  =  6'b110001;     //388pi/512
  assign cos2[388]  =  6'b111011;     //388pi/512
  assign sin2[389]  =  6'b110001;     //389pi/512
  assign cos2[389]  =  6'b111011;     //389pi/512
  assign sin2[390]  =  6'b110001;     //390pi/512
  assign cos2[390]  =  6'b111011;     //390pi/512
  assign sin2[391]  =  6'b110001;     //391pi/512
  assign cos2[391]  =  6'b111011;     //391pi/512
  assign sin2[392]  =  6'b110001;     //392pi/512
  assign cos2[392]  =  6'b111010;     //392pi/512
  assign sin2[393]  =  6'b110001;     //393pi/512
  assign cos2[393]  =  6'b111010;     //393pi/512
  assign sin2[394]  =  6'b110001;     //394pi/512
  assign cos2[394]  =  6'b111010;     //394pi/512
  assign sin2[395]  =  6'b110001;     //395pi/512
  assign cos2[395]  =  6'b111010;     //395pi/512
  assign sin2[396]  =  6'b110001;     //396pi/512
  assign cos2[396]  =  6'b111010;     //396pi/512
  assign sin2[397]  =  6'b110001;     //397pi/512
  assign cos2[397]  =  6'b111010;     //397pi/512
  assign sin2[398]  =  6'b110001;     //398pi/512
  assign cos2[398]  =  6'b111010;     //398pi/512
  assign sin2[399]  =  6'b110001;     //399pi/512
  assign cos2[399]  =  6'b111010;     //399pi/512
  assign sin2[400]  =  6'b110001;     //400pi/512
  assign cos2[400]  =  6'b111010;     //400pi/512
  assign sin2[401]  =  6'b110001;     //401pi/512
  assign cos2[401]  =  6'b111010;     //401pi/512
  assign sin2[402]  =  6'b110001;     //402pi/512
  assign cos2[402]  =  6'b111010;     //402pi/512
  assign sin2[403]  =  6'b110001;     //403pi/512
  assign cos2[403]  =  6'b111010;     //403pi/512
  assign sin2[404]  =  6'b110001;     //404pi/512
  assign cos2[404]  =  6'b111010;     //404pi/512
  assign sin2[405]  =  6'b110001;     //405pi/512
  assign cos2[405]  =  6'b111010;     //405pi/512
  assign sin2[406]  =  6'b110001;     //406pi/512
  assign cos2[406]  =  6'b111001;     //406pi/512
  assign sin2[407]  =  6'b110001;     //407pi/512
  assign cos2[407]  =  6'b111001;     //407pi/512
  assign sin2[408]  =  6'b110001;     //408pi/512
  assign cos2[408]  =  6'b111001;     //408pi/512
  assign sin2[409]  =  6'b110010;     //409pi/512
  assign cos2[409]  =  6'b111001;     //409pi/512
  assign sin2[410]  =  6'b110010;     //410pi/512
  assign cos2[410]  =  6'b111001;     //410pi/512
  assign sin2[411]  =  6'b110010;     //411pi/512
  assign cos2[411]  =  6'b111001;     //411pi/512
  assign sin2[412]  =  6'b110010;     //412pi/512
  assign cos2[412]  =  6'b111001;     //412pi/512
  assign sin2[413]  =  6'b110010;     //413pi/512
  assign cos2[413]  =  6'b111001;     //413pi/512
  assign sin2[414]  =  6'b110010;     //414pi/512
  assign cos2[414]  =  6'b111001;     //414pi/512
  assign sin2[415]  =  6'b110010;     //415pi/512
  assign cos2[415]  =  6'b111001;     //415pi/512
  assign sin2[416]  =  6'b110010;     //416pi/512
  assign cos2[416]  =  6'b111001;     //416pi/512
  assign sin2[417]  =  6'b110010;     //417pi/512
  assign cos2[417]  =  6'b111001;     //417pi/512
  assign sin2[418]  =  6'b110010;     //418pi/512
  assign cos2[418]  =  6'b111001;     //418pi/512
  assign sin2[419]  =  6'b110010;     //419pi/512
  assign cos2[419]  =  6'b111001;     //419pi/512
  assign sin2[420]  =  6'b110010;     //420pi/512
  assign cos2[420]  =  6'b111000;     //420pi/512
  assign sin2[421]  =  6'b110010;     //421pi/512
  assign cos2[421]  =  6'b111000;     //421pi/512
  assign sin2[422]  =  6'b110010;     //422pi/512
  assign cos2[422]  =  6'b111000;     //422pi/512
  assign sin2[423]  =  6'b110010;     //423pi/512
  assign cos2[423]  =  6'b111000;     //423pi/512
  assign sin2[424]  =  6'b110010;     //424pi/512
  assign cos2[424]  =  6'b111000;     //424pi/512
  assign sin2[425]  =  6'b110010;     //425pi/512
  assign cos2[425]  =  6'b111000;     //425pi/512
  assign sin2[426]  =  6'b110010;     //426pi/512
  assign cos2[426]  =  6'b111000;     //426pi/512
  assign sin2[427]  =  6'b110010;     //427pi/512
  assign cos2[427]  =  6'b111000;     //427pi/512
  assign sin2[428]  =  6'b110010;     //428pi/512
  assign cos2[428]  =  6'b111000;     //428pi/512
  assign sin2[429]  =  6'b110010;     //429pi/512
  assign cos2[429]  =  6'b111000;     //429pi/512
  assign sin2[430]  =  6'b110010;     //430pi/512
  assign cos2[430]  =  6'b111000;     //430pi/512
  assign sin2[431]  =  6'b110010;     //431pi/512
  assign cos2[431]  =  6'b111000;     //431pi/512
  assign sin2[432]  =  6'b110010;     //432pi/512
  assign cos2[432]  =  6'b111000;     //432pi/512
  assign sin2[433]  =  6'b110010;     //433pi/512
  assign cos2[433]  =  6'b111000;     //433pi/512
  assign sin2[434]  =  6'b110010;     //434pi/512
  assign cos2[434]  =  6'b111000;     //434pi/512
  assign sin2[435]  =  6'b110010;     //435pi/512
  assign cos2[435]  =  6'b110111;     //435pi/512
  assign sin2[436]  =  6'b110011;     //436pi/512
  assign cos2[436]  =  6'b110111;     //436pi/512
  assign sin2[437]  =  6'b110011;     //437pi/512
  assign cos2[437]  =  6'b110111;     //437pi/512
  assign sin2[438]  =  6'b110011;     //438pi/512
  assign cos2[438]  =  6'b110111;     //438pi/512
  assign sin2[439]  =  6'b110011;     //439pi/512
  assign cos2[439]  =  6'b110111;     //439pi/512
  assign sin2[440]  =  6'b110011;     //440pi/512
  assign cos2[440]  =  6'b110111;     //440pi/512
  assign sin2[441]  =  6'b110011;     //441pi/512
  assign cos2[441]  =  6'b110111;     //441pi/512
  assign sin2[442]  =  6'b110011;     //442pi/512
  assign cos2[442]  =  6'b110111;     //442pi/512
  assign sin2[443]  =  6'b110011;     //443pi/512
  assign cos2[443]  =  6'b110111;     //443pi/512
  assign sin2[444]  =  6'b110011;     //444pi/512
  assign cos2[444]  =  6'b110111;     //444pi/512
  assign sin2[445]  =  6'b110011;     //445pi/512
  assign cos2[445]  =  6'b110111;     //445pi/512
  assign sin2[446]  =  6'b110011;     //446pi/512
  assign cos2[446]  =  6'b110111;     //446pi/512
  assign sin2[447]  =  6'b110011;     //447pi/512
  assign cos2[447]  =  6'b110111;     //447pi/512
  assign sin2[448]  =  6'b110011;     //448pi/512
  assign cos2[448]  =  6'b110111;     //448pi/512
  assign sin2[449]  =  6'b110011;     //449pi/512
  assign cos2[449]  =  6'b110111;     //449pi/512
  assign sin2[450]  =  6'b110011;     //450pi/512
  assign cos2[450]  =  6'b110110;     //450pi/512
  assign sin2[451]  =  6'b110011;     //451pi/512
  assign cos2[451]  =  6'b110110;     //451pi/512
  assign sin2[452]  =  6'b110011;     //452pi/512
  assign cos2[452]  =  6'b110110;     //452pi/512
  assign sin2[453]  =  6'b110011;     //453pi/512
  assign cos2[453]  =  6'b110110;     //453pi/512
  assign sin2[454]  =  6'b110011;     //454pi/512
  assign cos2[454]  =  6'b110110;     //454pi/512
  assign sin2[455]  =  6'b110011;     //455pi/512
  assign cos2[455]  =  6'b110110;     //455pi/512
  assign sin2[456]  =  6'b110011;     //456pi/512
  assign cos2[456]  =  6'b110110;     //456pi/512
  assign sin2[457]  =  6'b110011;     //457pi/512
  assign cos2[457]  =  6'b110110;     //457pi/512
  assign sin2[458]  =  6'b110100;     //458pi/512
  assign cos2[458]  =  6'b110110;     //458pi/512
  assign sin2[459]  =  6'b110100;     //459pi/512
  assign cos2[459]  =  6'b110110;     //459pi/512
  assign sin2[460]  =  6'b110100;     //460pi/512
  assign cos2[460]  =  6'b110110;     //460pi/512
  assign sin2[461]  =  6'b110100;     //461pi/512
  assign cos2[461]  =  6'b110110;     //461pi/512
  assign sin2[462]  =  6'b110100;     //462pi/512
  assign cos2[462]  =  6'b110110;     //462pi/512
  assign sin2[463]  =  6'b110100;     //463pi/512
  assign cos2[463]  =  6'b110110;     //463pi/512
  assign sin2[464]  =  6'b110100;     //464pi/512
  assign cos2[464]  =  6'b110110;     //464pi/512
  assign sin2[465]  =  6'b110100;     //465pi/512
  assign cos2[465]  =  6'b110110;     //465pi/512
  assign sin2[466]  =  6'b110100;     //466pi/512
  assign cos2[466]  =  6'b110101;     //466pi/512
  assign sin2[467]  =  6'b110100;     //467pi/512
  assign cos2[467]  =  6'b110101;     //467pi/512
  assign sin2[468]  =  6'b110100;     //468pi/512
  assign cos2[468]  =  6'b110101;     //468pi/512
  assign sin2[469]  =  6'b110100;     //469pi/512
  assign cos2[469]  =  6'b110101;     //469pi/512
  assign sin2[470]  =  6'b110100;     //470pi/512
  assign cos2[470]  =  6'b110101;     //470pi/512
  assign sin2[471]  =  6'b110100;     //471pi/512
  assign cos2[471]  =  6'b110101;     //471pi/512
  assign sin2[472]  =  6'b110100;     //472pi/512
  assign cos2[472]  =  6'b110101;     //472pi/512
  assign sin2[473]  =  6'b110100;     //473pi/512
  assign cos2[473]  =  6'b110101;     //473pi/512
  assign sin2[474]  =  6'b110100;     //474pi/512
  assign cos2[474]  =  6'b110101;     //474pi/512
  assign sin2[475]  =  6'b110100;     //475pi/512
  assign cos2[475]  =  6'b110101;     //475pi/512
  assign sin2[476]  =  6'b110100;     //476pi/512
  assign cos2[476]  =  6'b110101;     //476pi/512
  assign sin2[477]  =  6'b110101;     //477pi/512
  assign cos2[477]  =  6'b110101;     //477pi/512
  assign sin2[478]  =  6'b110101;     //478pi/512
  assign cos2[478]  =  6'b110101;     //478pi/512
  assign sin2[479]  =  6'b110101;     //479pi/512
  assign cos2[479]  =  6'b110101;     //479pi/512
  assign sin2[480]  =  6'b110101;     //480pi/512
  assign cos2[480]  =  6'b110101;     //480pi/512
  assign sin2[481]  =  6'b110101;     //481pi/512
  assign cos2[481]  =  6'b110101;     //481pi/512
  assign sin2[482]  =  6'b110101;     //482pi/512
  assign cos2[482]  =  6'b110101;     //482pi/512
  assign sin2[483]  =  6'b110101;     //483pi/512
  assign cos2[483]  =  6'b110101;     //483pi/512
  assign sin2[484]  =  6'b110101;     //484pi/512
  assign cos2[484]  =  6'b110100;     //484pi/512
  assign sin2[485]  =  6'b110101;     //485pi/512
  assign cos2[485]  =  6'b110100;     //485pi/512
  assign sin2[486]  =  6'b110101;     //486pi/512
  assign cos2[486]  =  6'b110100;     //486pi/512
  assign sin2[487]  =  6'b110101;     //487pi/512
  assign cos2[487]  =  6'b110100;     //487pi/512
  assign sin2[488]  =  6'b110101;     //488pi/512
  assign cos2[488]  =  6'b110100;     //488pi/512
  assign sin2[489]  =  6'b110101;     //489pi/512
  assign cos2[489]  =  6'b110100;     //489pi/512
  assign sin2[490]  =  6'b110101;     //490pi/512
  assign cos2[490]  =  6'b110100;     //490pi/512
  assign sin2[491]  =  6'b110101;     //491pi/512
  assign cos2[491]  =  6'b110100;     //491pi/512
  assign sin2[492]  =  6'b110101;     //492pi/512
  assign cos2[492]  =  6'b110100;     //492pi/512
  assign sin2[493]  =  6'b110101;     //493pi/512
  assign cos2[493]  =  6'b110100;     //493pi/512
  assign sin2[494]  =  6'b110101;     //494pi/512
  assign cos2[494]  =  6'b110100;     //494pi/512
  assign sin2[495]  =  6'b110110;     //495pi/512
  assign cos2[495]  =  6'b110100;     //495pi/512
  assign sin2[496]  =  6'b110110;     //496pi/512
  assign cos2[496]  =  6'b110100;     //496pi/512
  assign sin2[497]  =  6'b110110;     //497pi/512
  assign cos2[497]  =  6'b110100;     //497pi/512
  assign sin2[498]  =  6'b110110;     //498pi/512
  assign cos2[498]  =  6'b110100;     //498pi/512
  assign sin2[499]  =  6'b110110;     //499pi/512
  assign cos2[499]  =  6'b110100;     //499pi/512
  assign sin2[500]  =  6'b110110;     //500pi/512
  assign cos2[500]  =  6'b110100;     //500pi/512
  assign sin2[501]  =  6'b110110;     //501pi/512
  assign cos2[501]  =  6'b110100;     //501pi/512
  assign sin2[502]  =  6'b110110;     //502pi/512
  assign cos2[502]  =  6'b110100;     //502pi/512
  assign sin2[503]  =  6'b110110;     //503pi/512
  assign cos2[503]  =  6'b110011;     //503pi/512
  assign sin2[504]  =  6'b110110;     //504pi/512
  assign cos2[504]  =  6'b110011;     //504pi/512
  assign sin2[505]  =  6'b110110;     //505pi/512
  assign cos2[505]  =  6'b110011;     //505pi/512
  assign sin2[506]  =  6'b110110;     //506pi/512
  assign cos2[506]  =  6'b110011;     //506pi/512
  assign sin2[507]  =  6'b110110;     //507pi/512
  assign cos2[507]  =  6'b110011;     //507pi/512
  assign sin2[508]  =  6'b110110;     //508pi/512
  assign cos2[508]  =  6'b110011;     //508pi/512
  assign sin2[509]  =  6'b110110;     //509pi/512
  assign cos2[509]  =  6'b110011;     //509pi/512
  assign sin2[510]  =  6'b110110;     //510pi/512
  assign cos2[510]  =  6'b110011;     //510pi/512
  assign sin2[511]  =  6'b110111;     //511pi/512
  assign cos2[511]  =  6'b110011;     //511pi/512
 
endmodule