
module modifying_adder
	#(parameter bit_width=16, SIZE = 4)(
    input   [3:0] stage_FFT,
    
    input   signed [bit_width-1:0] xin1,
    input   signed [bit_width-1:0] yin1,
	input   signed [bit_width-1:0] xin2,
	input   signed [bit_width-1:0] yin2,
    input   signed [bit_width-1:0] xin3,
	input   signed [bit_width-1:0] yin3,
    input   en,
    input   delay,

    output  signed [bit_width-1:0]  xout1,
	output  signed [bit_width-1:0]  yout1,
    output  signed [bit_width-1:0]  xout2,
	output  signed [bit_width-1:0]  yout2
    
   );
   
  assign xout1 = (en || delay)?  xin1 + xin2 : xout1;
  assign yout1 = (en || delay)?  yin1 + yin2 : yout1;
 // assign xout2 = (stage_FFT == SIZE && en)? xin1 + xin3  : en?  xin1-xin2  :xout2;
 // assign yout2 = (stage_FFT == SIZE && en)? yin1 + yin3  : en?  yin1-yin2  :yout2;
  
  assign xout2 = (stage_FFT >= SIZE && (en || delay))? xin1 + xin3  : (en || delay)? xin1-xin2 : xout2 ;
  assign yout2 = (stage_FFT >= SIZE && (en || delay))? yin1 + yin3  : (en || delay)? yin1-yin2 : yout2 ; 

endmodule