module  tw_factor_for_8th #(parameter stage_FFT = 2, SIZE =10, word_length_tw = 14) (
    input            clk,
    input            en_rd, 
    input   [stage_FFT-2:0]   rd_ptr_angle,

    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );


reg signed [word_length_tw-1:0]  cos  [127:0];
reg signed [word_length_tw-1:0]  sin  [127:0];


//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd  ) begin
                  cos_data           <= cos   [rd_ptr_angle];
                  sin_data           <= sin   [rd_ptr_angle];
             end 
        end

//--------------------------------handle read tw factor------------------------------

initial begin
   sin[0]  =  14'b00000000000000;     //0pi/1024
   cos[0]  =  14'b01000000000000;     //0pi/1024
   sin[1]  =  14'b11111110011011;     //8pi/1024
   cos[1]  =  14'b00111111111110;     //8pi/1024
   sin[2]  =  14'b11111100110111;     //16pi/1024
   cos[2]  =  14'b00111111111011;     //16pi/1024
   sin[3]  =  14'b11111011010011;     //24pi/1024
   cos[3]  =  14'b00111111110100;     //24pi/1024
   sin[4]  =  14'b11111001101111;     //32pi/1024
   cos[4]  =  14'b00111111101100;     //32pi/1024
   sin[5]  =  14'b11111000001011;     //40pi/1024
   cos[5]  =  14'b00111111100001;     //40pi/1024
   sin[6]  =  14'b11110110100111;     //48pi/1024
   cos[6]  =  14'b00111111010011;     //48pi/1024
   sin[7]  =  14'b11110101000100;     //56pi/1024
   cos[7]  =  14'b00111111000011;     //56pi/1024
   sin[8]  =  14'b11110011100001;     //64pi/1024
   cos[8]  =  14'b00111110110001;     //64pi/1024
   sin[9]  =  14'b11110001111111;     //72pi/1024
   cos[9]  =  14'b00111110011100;     //72pi/1024
   sin[10]  =  14'b11110000011101;     //80pi/1024
   cos[10]  =  14'b00111110000101;     //80pi/1024
   sin[11]  =  14'b11101110111100;     //88pi/1024
   cos[11]  =  14'b00111101101011;     //88pi/1024
   sin[12]  =  14'b11101101011011;     //96pi/1024
   cos[12]  =  14'b00111101001111;     //96pi/1024
   sin[13]  =  14'b11101011111011;     //104pi/1024
   cos[13]  =  14'b00111100110001;     //104pi/1024
   sin[14]  =  14'b11101010011100;     //112pi/1024
   cos[14]  =  14'b00111100010000;     //112pi/1024
   sin[15]  =  14'b11101000111110;     //120pi/1024
   cos[15]  =  14'b00111011101101;     //120pi/1024
   sin[16]  =  14'b11100111100001;     //128pi/1024
   cos[16]  =  14'b00111011001000;     //128pi/1024
   sin[17]  =  14'b11100110000100;     //136pi/1024
   cos[17]  =  14'b00111010100000;     //136pi/1024
   sin[18]  =  14'b11100100101001;     //144pi/1024
   cos[18]  =  14'b00111001110110;     //144pi/1024
   sin[19]  =  14'b11100011001110;     //152pi/1024
   cos[19]  =  14'b00111001001010;     //152pi/1024
   sin[20]  =  14'b11100001110101;     //160pi/1024
   cos[20]  =  14'b00111000011100;     //160pi/1024
   sin[21]  =  14'b11100000011101;     //168pi/1024
   cos[21]  =  14'b00110111101011;     //168pi/1024
   sin[22]  =  14'b11011111000110;     //176pi/1024
   cos[22]  =  14'b00110110111001;     //176pi/1024
   sin[23]  =  14'b11011101110001;     //184pi/1024
   cos[23]  =  14'b00110110000100;     //184pi/1024
   sin[24]  =  14'b11011100011100;     //192pi/1024
   cos[24]  =  14'b00110101001101;     //192pi/1024
   sin[25]  =  14'b11011011001001;     //200pi/1024
   cos[25]  =  14'b00110100010100;     //200pi/1024
   sin[26]  =  14'b11011001111000;     //208pi/1024
   cos[26]  =  14'b00110011011001;     //208pi/1024
   sin[27]  =  14'b11011000101000;     //216pi/1024
   cos[27]  =  14'b00110010011101;     //216pi/1024
   sin[28]  =  14'b11010111011010;     //224pi/1024
   cos[28]  =  14'b00110001011110;     //224pi/1024
   sin[29]  =  14'b11010110001101;     //232pi/1024
   cos[29]  =  14'b00110000011101;     //232pi/1024
   sin[30]  =  14'b11010101000001;     //240pi/1024
   cos[30]  =  14'b00101111011010;     //240pi/1024
   sin[31]  =  14'b11010011111000;     //248pi/1024
   cos[31]  =  14'b00101110010110;     //248pi/1024
   sin[32]  =  14'b11010010110000;     //256pi/1024
   cos[32]  =  14'b00101101010000;     //256pi/1024
   sin[33]  =  14'b11010001101001;     //264pi/1024
   cos[33]  =  14'b00101100001000;     //264pi/1024
   sin[34]  =  14'b11010000100101;     //272pi/1024
   cos[34]  =  14'b00101010111110;     //272pi/1024
   sin[35]  =  14'b11001111100010;     //280pi/1024
   cos[35]  =  14'b00101001110011;     //280pi/1024
   sin[36]  =  14'b11001110100010;     //288pi/1024
   cos[36]  =  14'b00101000100110;     //288pi/1024
   sin[37]  =  14'b11001101100011;     //296pi/1024
   cos[37]  =  14'b00100111010111;     //296pi/1024
   sin[38]  =  14'b11001100100110;     //304pi/1024
   cos[38]  =  14'b00100110000111;     //304pi/1024
   sin[39]  =  14'b11001011101011;     //312pi/1024
   cos[39]  =  14'b00100100110110;     //312pi/1024
   sin[40]  =  14'b11001010110010;     //320pi/1024
   cos[40]  =  14'b00100011100011;     //320pi/1024
   sin[41]  =  14'b11001001111011;     //328pi/1024
   cos[41]  =  14'b00100010001111;     //328pi/1024
   sin[42]  =  14'b11001001000111;     //336pi/1024
   cos[42]  =  14'b00100000111001;     //336pi/1024
   sin[43]  =  14'b11001000010100;     //344pi/1024
   cos[43]  =  14'b00011111100010;     //344pi/1024
   sin[44]  =  14'b11000111100100;     //352pi/1024
   cos[44]  =  14'b00011110001010;     //352pi/1024
   sin[45]  =  14'b11000110110101;     //360pi/1024
   cos[45]  =  14'b00011100110001;     //360pi/1024
   sin[46]  =  14'b11000110001001;     //368pi/1024
   cos[46]  =  14'b00011011010111;     //368pi/1024
   sin[47]  =  14'b11000101011111;     //376pi/1024
   cos[47]  =  14'b00011001111011;     //376pi/1024
   sin[48]  =  14'b11000100111000;     //384pi/1024
   cos[48]  =  14'b00011000011111;     //384pi/1024
   sin[49]  =  14'b11000100010010;     //392pi/1024
   cos[49]  =  14'b00010111000010;     //392pi/1024
   sin[50]  =  14'b11000011101111;     //400pi/1024
   cos[50]  =  14'b00010101100011;     //400pi/1024
   sin[51]  =  14'b11000011001111;     //408pi/1024
   cos[51]  =  14'b00010100000100;     //408pi/1024
   sin[52]  =  14'b11000010110000;     //416pi/1024
   cos[52]  =  14'b00010010100101;     //416pi/1024
   sin[53]  =  14'b11000010010100;     //424pi/1024
   cos[53]  =  14'b00010001000100;     //424pi/1024
   sin[54]  =  14'b11000001111011;     //432pi/1024
   cos[54]  =  14'b00001111100011;     //432pi/1024
   sin[55]  =  14'b11000001100100;     //440pi/1024
   cos[55]  =  14'b00001110000001;     //440pi/1024
   sin[56]  =  14'b11000001001111;     //448pi/1024
   cos[56]  =  14'b00001100011111;     //448pi/1024
   sin[57]  =  14'b11000000111100;     //456pi/1024
   cos[57]  =  14'b00001010111100;     //456pi/1024
   sin[58]  =  14'b11000000101100;     //464pi/1024
   cos[58]  =  14'b00001001011001;     //464pi/1024
   sin[59]  =  14'b11000000011111;     //472pi/1024
   cos[59]  =  14'b00000111110101;     //472pi/1024
   sin[60]  =  14'b11000000010100;     //480pi/1024
   cos[60]  =  14'b00000110010001;     //480pi/1024
   sin[61]  =  14'b11000000001011;     //488pi/1024
   cos[61]  =  14'b00000100101101;     //488pi/1024
   sin[62]  =  14'b11000000000101;     //496pi/1024
   cos[62]  =  14'b00000011001000;     //496pi/1024
   sin[63]  =  14'b11000000000001;     //504pi/1024
   cos[63]  =  14'b00000001100100;     //504pi/1024
   sin[64]  =  14'b11000000000000;     //512pi/1024
   cos[64]  =  14'b00000000000000;     //512pi/1024
   sin[65]  =  14'b11000000000001;     //520pi/1024
   cos[65]  =  14'b11111110011011;     //520pi/1024
   sin[66]  =  14'b11000000000101;     //528pi/1024
   cos[66]  =  14'b11111100110111;     //528pi/1024
   sin[67]  =  14'b11000000001011;     //536pi/1024
   cos[67]  =  14'b11111011010011;     //536pi/1024
   sin[68]  =  14'b11000000010100;     //544pi/1024
   cos[68]  =  14'b11111001101111;     //544pi/1024
   sin[69]  =  14'b11000000011111;     //552pi/1024
   cos[69]  =  14'b11111000001011;     //552pi/1024
   sin[70]  =  14'b11000000101100;     //560pi/1024
   cos[70]  =  14'b11110110100111;     //560pi/1024
   sin[71]  =  14'b11000000111100;     //568pi/1024
   cos[71]  =  14'b11110101000100;     //568pi/1024
   sin[72]  =  14'b11000001001111;     //576pi/1024
   cos[72]  =  14'b11110011100001;     //576pi/1024
   sin[73]  =  14'b11000001100100;     //584pi/1024
   cos[73]  =  14'b11110001111111;     //584pi/1024
   sin[74]  =  14'b11000001111011;     //592pi/1024
   cos[74]  =  14'b11110000011101;     //592pi/1024
   sin[75]  =  14'b11000010010100;     //600pi/1024
   cos[75]  =  14'b11101110111100;     //600pi/1024
   sin[76]  =  14'b11000010110000;     //608pi/1024
   cos[76]  =  14'b11101101011011;     //608pi/1024
   sin[77]  =  14'b11000011001111;     //616pi/1024
   cos[77]  =  14'b11101011111011;     //616pi/1024
   sin[78]  =  14'b11000011101111;     //624pi/1024
   cos[78]  =  14'b11101010011100;     //624pi/1024
   sin[79]  =  14'b11000100010010;     //632pi/1024
   cos[79]  =  14'b11101000111110;     //632pi/1024
   sin[80]  =  14'b11000100111000;     //640pi/1024
   cos[80]  =  14'b11100111100001;     //640pi/1024
   sin[81]  =  14'b11000101011111;     //648pi/1024
   cos[81]  =  14'b11100110000100;     //648pi/1024
   sin[82]  =  14'b11000110001001;     //656pi/1024
   cos[82]  =  14'b11100100101001;     //656pi/1024
   sin[83]  =  14'b11000110110101;     //664pi/1024
   cos[83]  =  14'b11100011001110;     //664pi/1024
   sin[84]  =  14'b11000111100100;     //672pi/1024
   cos[84]  =  14'b11100001110101;     //672pi/1024
   sin[85]  =  14'b11001000010100;     //680pi/1024
   cos[85]  =  14'b11100000011101;     //680pi/1024
   sin[86]  =  14'b11001001000111;     //688pi/1024
   cos[86]  =  14'b11011111000110;     //688pi/1024
   sin[87]  =  14'b11001001111011;     //696pi/1024
   cos[87]  =  14'b11011101110001;     //696pi/1024
   sin[88]  =  14'b11001010110010;     //704pi/1024
   cos[88]  =  14'b11011100011100;     //704pi/1024
   sin[89]  =  14'b11001011101011;     //712pi/1024
   cos[89]  =  14'b11011011001001;     //712pi/1024
   sin[90]  =  14'b11001100100110;     //720pi/1024
   cos[90]  =  14'b11011001111000;     //720pi/1024
   sin[91]  =  14'b11001101100011;     //728pi/1024
   cos[91]  =  14'b11011000101000;     //728pi/1024
   sin[92]  =  14'b11001110100010;     //736pi/1024
   cos[92]  =  14'b11010111011010;     //736pi/1024
   sin[93]  =  14'b11001111100010;     //744pi/1024
   cos[93]  =  14'b11010110001101;     //744pi/1024
   sin[94]  =  14'b11010000100101;     //752pi/1024
   cos[94]  =  14'b11010101000001;     //752pi/1024
   sin[95]  =  14'b11010001101001;     //760pi/1024
   cos[95]  =  14'b11010011111000;     //760pi/1024
   sin[96]  =  14'b11010010110000;     //768pi/1024
   cos[96]  =  14'b11010010110000;     //768pi/1024
   sin[97]  =  14'b11010011111000;     //776pi/1024
   cos[97]  =  14'b11010001101001;     //776pi/1024
   sin[98]  =  14'b11010101000001;     //784pi/1024
   cos[98]  =  14'b11010000100101;     //784pi/1024
   sin[99]  =  14'b11010110001101;     //792pi/1024
   cos[99]  =  14'b11001111100010;     //792pi/1024
   sin[100]  =  14'b11010111011010;     //800pi/1024
   cos[100]  =  14'b11001110100010;     //800pi/1024
   sin[101]  =  14'b11011000101000;     //808pi/1024
   cos[101]  =  14'b11001101100011;     //808pi/1024
   sin[102]  =  14'b11011001111000;     //816pi/1024
   cos[102]  =  14'b11001100100110;     //816pi/1024
   sin[103]  =  14'b11011011001001;     //824pi/1024
   cos[103]  =  14'b11001011101011;     //824pi/1024
   sin[104]  =  14'b11011100011100;     //832pi/1024
   cos[104]  =  14'b11001010110010;     //832pi/1024
   sin[105]  =  14'b11011101110001;     //840pi/1024
   cos[105]  =  14'b11001001111011;     //840pi/1024
   sin[106]  =  14'b11011111000110;     //848pi/1024
   cos[106]  =  14'b11001001000111;     //848pi/1024
   sin[107]  =  14'b11100000011101;     //856pi/1024
   cos[107]  =  14'b11001000010100;     //856pi/1024
   sin[108]  =  14'b11100001110101;     //864pi/1024
   cos[108]  =  14'b11000111100100;     //864pi/1024
   sin[109]  =  14'b11100011001110;     //872pi/1024
   cos[109]  =  14'b11000110110101;     //872pi/1024
   sin[110]  =  14'b11100100101001;     //880pi/1024
   cos[110]  =  14'b11000110001001;     //880pi/1024
   sin[111]  =  14'b11100110000100;     //888pi/1024
   cos[111]  =  14'b11000101011111;     //888pi/1024
   sin[112]  =  14'b11100111100001;     //896pi/1024
   cos[112]  =  14'b11000100111000;     //896pi/1024
   sin[113]  =  14'b11101000111110;     //904pi/1024
   cos[113]  =  14'b11000100010010;     //904pi/1024
   sin[114]  =  14'b11101010011100;     //912pi/1024
   cos[114]  =  14'b11000011101111;     //912pi/1024
   sin[115]  =  14'b11101011111011;     //920pi/1024
   cos[115]  =  14'b11000011001111;     //920pi/1024
   sin[116]  =  14'b11101101011011;     //928pi/1024
   cos[116]  =  14'b11000010110000;     //928pi/1024
   sin[117]  =  14'b11101110111100;     //936pi/1024
   cos[117]  =  14'b11000010010100;     //936pi/1024
   sin[118]  =  14'b11110000011101;     //944pi/1024
   cos[118]  =  14'b11000001111011;     //944pi/1024
   sin[119]  =  14'b11110001111111;     //952pi/1024
   cos[119]  =  14'b11000001100100;     //952pi/1024
   sin[120]  =  14'b11110011100001;     //960pi/1024
   cos[120]  =  14'b11000001001111;     //960pi/1024
   sin[121]  =  14'b11110101000100;     //968pi/1024
   cos[121]  =  14'b11000000111100;     //968pi/1024
   sin[122]  =  14'b11110110100111;     //976pi/1024
   cos[122]  =  14'b11000000101100;     //976pi/1024
   sin[123]  =  14'b11111000001011;     //984pi/1024
   cos[123]  =  14'b11000000011111;     //984pi/1024
   sin[124]  =  14'b11111001101111;     //992pi/1024
   cos[124]  =  14'b11000000010100;     //992pi/1024
   sin[125]  =  14'b11111011010011;     //1000pi/1024
   cos[125]  =  14'b11000000001011;     //1000pi/1024
   sin[126]  =  14'b11111100110111;     //1008pi/1024
   cos[126]  =  14'b11000000000101;     //1008pi/1024
   sin[127]  =  14'b11111110011011;     //1016pi/1024
   cos[127]  =  14'b11000000000001;     //1016pi/1024
end
endmodule