module  M_TWIDLE_14_bit #(parameter SIZE =10) (
    input            clk,
    input            en, 
    input   [10:0]   rd_ptr_angle,

    output  reg signed [13:0]   cos_data,
    output  reg signed [13:0]   sin_data
 );


reg signed [13:0]  cos  [1023:0];
reg signed [13:0]  sin  [1023:0];

wire  en_rd;

wire       [10:0]  rd_ptr;

shift_register # ( .width (11), .depth (2)) shift_register1(
         .clk(clk),
         .rst_n(rst_n), 
         .in_data(rd_ptr_angle),
         .out_data(rd_ptr)
);
shift_register # ( .width (1), .depth (2)) shift_register2(
         .clk(clk),
         .rst_n(rst_n), 
         .in_data(en),
         .out_data(en_rd)
);
always @(posedge clk ) begin
  if (en_rd) begin
    cos_data <=   cos [rd_ptr];
    sin_data <=   sin [rd_ptr];
  end 
end

initial begin
   sin[0]  =  14'b00000000000000;     //0pi/512
   cos[0]  =  14'b01000000000000;     //0pi/512
   sin[1]  =  14'b11111111100111;     //1pi/512
   cos[1]  =  14'b00111111111111;     //1pi/512
   sin[2]  =  14'b11111111001110;     //2pi/512
   cos[2]  =  14'b00111111111111;     //2pi/512
   sin[3]  =  14'b11111110110101;     //3pi/512
   cos[3]  =  14'b00111111111111;     //3pi/512
   sin[4]  =  14'b11111110011011;     //4pi/512
   cos[4]  =  14'b00111111111110;     //4pi/512
   sin[5]  =  14'b11111110000010;     //5pi/512
   cos[5]  =  14'b00111111111110;     //5pi/512
   sin[6]  =  14'b11111101101001;     //6pi/512
   cos[6]  =  14'b00111111111101;     //6pi/512
   sin[7]  =  14'b11111101010000;     //7pi/512
   cos[7]  =  14'b00111111111100;     //7pi/512
   sin[8]  =  14'b11111100110111;     //8pi/512
   cos[8]  =  14'b00111111111011;     //8pi/512
   sin[9]  =  14'b11111100011110;     //9pi/512
   cos[9]  =  14'b00111111111001;     //9pi/512
   sin[10]  =  14'b11111100000101;     //10pi/512
   cos[10]  =  14'b00111111111000;     //10pi/512
   sin[11]  =  14'b11111011101100;     //11pi/512
   cos[11]  =  14'b00111111110110;     //11pi/512
   sin[12]  =  14'b11111011010011;     //12pi/512
   cos[12]  =  14'b00111111110100;     //12pi/512
   sin[13]  =  14'b11111010111010;     //13pi/512
   cos[13]  =  14'b00111111110010;     //13pi/512
   sin[14]  =  14'b11111010100001;     //14pi/512
   cos[14]  =  14'b00111111110000;     //14pi/512
   sin[15]  =  14'b11111010001000;     //15pi/512
   cos[15]  =  14'b00111111101110;     //15pi/512
   sin[16]  =  14'b11111001101111;     //16pi/512
   cos[16]  =  14'b00111111101100;     //16pi/512
   sin[17]  =  14'b11111001010110;     //17pi/512
   cos[17]  =  14'b00111111101001;     //17pi/512
   sin[18]  =  14'b11111000111101;     //18pi/512
   cos[18]  =  14'b00111111100111;     //18pi/512
   sin[19]  =  14'b11111000100100;     //19pi/512
   cos[19]  =  14'b00111111100100;     //19pi/512
   sin[20]  =  14'b11111000001011;     //20pi/512
   cos[20]  =  14'b00111111100001;     //20pi/512
   sin[21]  =  14'b11110111110010;     //21pi/512
   cos[21]  =  14'b00111111011110;     //21pi/512
   sin[22]  =  14'b11110111011001;     //22pi/512
   cos[22]  =  14'b00111111011010;     //22pi/512
   sin[23]  =  14'b11110111000000;     //23pi/512
   cos[23]  =  14'b00111111010111;     //23pi/512
   sin[24]  =  14'b11110110100111;     //24pi/512
   cos[24]  =  14'b00111111010011;     //24pi/512
   sin[25]  =  14'b11110110001110;     //25pi/512
   cos[25]  =  14'b00111111001111;     //25pi/512
   sin[26]  =  14'b11110101110101;     //26pi/512
   cos[26]  =  14'b00111111001011;     //26pi/512
   sin[27]  =  14'b11110101011101;     //27pi/512
   cos[27]  =  14'b00111111000111;     //27pi/512
   sin[28]  =  14'b11110101000100;     //28pi/512
   cos[28]  =  14'b00111111000011;     //28pi/512
   sin[29]  =  14'b11110100101011;     //29pi/512
   cos[29]  =  14'b00111110111111;     //29pi/512
   sin[30]  =  14'b11110100010010;     //30pi/512
   cos[30]  =  14'b00111110111010;     //30pi/512
   sin[31]  =  14'b11110011111010;     //31pi/512
   cos[31]  =  14'b00111110110110;     //31pi/512
   sin[32]  =  14'b11110011100001;     //32pi/512
   cos[32]  =  14'b00111110110001;     //32pi/512
   sin[33]  =  14'b11110011001000;     //33pi/512
   cos[33]  =  14'b00111110101100;     //33pi/512
   sin[34]  =  14'b11110010110000;     //34pi/512
   cos[34]  =  14'b00111110100111;     //34pi/512
   sin[35]  =  14'b11110010010111;     //35pi/512
   cos[35]  =  14'b00111110100001;     //35pi/512
   sin[36]  =  14'b11110001111111;     //36pi/512
   cos[36]  =  14'b00111110011100;     //36pi/512
   sin[37]  =  14'b11110001100110;     //37pi/512
   cos[37]  =  14'b00111110010110;     //37pi/512
   sin[38]  =  14'b11110001001110;     //38pi/512
   cos[38]  =  14'b00111110010001;     //38pi/512
   sin[39]  =  14'b11110000110101;     //39pi/512
   cos[39]  =  14'b00111110001011;     //39pi/512
   sin[40]  =  14'b11110000011101;     //40pi/512
   cos[40]  =  14'b00111110000101;     //40pi/512
   sin[41]  =  14'b11110000000100;     //41pi/512
   cos[41]  =  14'b00111101111111;     //41pi/512
   sin[42]  =  14'b11101111101100;     //42pi/512
   cos[42]  =  14'b00111101111000;     //42pi/512
   sin[43]  =  14'b11101111010100;     //43pi/512
   cos[43]  =  14'b00111101110010;     //43pi/512
   sin[44]  =  14'b11101110111100;     //44pi/512
   cos[44]  =  14'b00111101101011;     //44pi/512
   sin[45]  =  14'b11101110100011;     //45pi/512
   cos[45]  =  14'b00111101100100;     //45pi/512
   sin[46]  =  14'b11101110001011;     //46pi/512
   cos[46]  =  14'b00111101011101;     //46pi/512
   sin[47]  =  14'b11101101110011;     //47pi/512
   cos[47]  =  14'b00111101010110;     //47pi/512
   sin[48]  =  14'b11101101011011;     //48pi/512
   cos[48]  =  14'b00111101001111;     //48pi/512
   sin[49]  =  14'b11101101000011;     //49pi/512
   cos[49]  =  14'b00111101001000;     //49pi/512
   sin[50]  =  14'b11101100101011;     //50pi/512
   cos[50]  =  14'b00111101000000;     //50pi/512
   sin[51]  =  14'b11101100010011;     //51pi/512
   cos[51]  =  14'b00111100111001;     //51pi/512
   sin[52]  =  14'b11101011111011;     //52pi/512
   cos[52]  =  14'b00111100110001;     //52pi/512
   sin[53]  =  14'b11101011100011;     //53pi/512
   cos[53]  =  14'b00111100101001;     //53pi/512
   sin[54]  =  14'b11101011001100;     //54pi/512
   cos[54]  =  14'b00111100100001;     //54pi/512
   sin[55]  =  14'b11101010110100;     //55pi/512
   cos[55]  =  14'b00111100011000;     //55pi/512
   sin[56]  =  14'b11101010011100;     //56pi/512
   cos[56]  =  14'b00111100010000;     //56pi/512
   sin[57]  =  14'b11101010000100;     //57pi/512
   cos[57]  =  14'b00111100001000;     //57pi/512
   sin[58]  =  14'b11101001101101;     //58pi/512
   cos[58]  =  14'b00111011111111;     //58pi/512
   sin[59]  =  14'b11101001010101;     //59pi/512
   cos[59]  =  14'b00111011110110;     //59pi/512
   sin[60]  =  14'b11101000111110;     //60pi/512
   cos[60]  =  14'b00111011101101;     //60pi/512
   sin[61]  =  14'b11101000100110;     //61pi/512
   cos[61]  =  14'b00111011100100;     //61pi/512
   sin[62]  =  14'b11101000001111;     //62pi/512
   cos[62]  =  14'b00111011011011;     //62pi/512
   sin[63]  =  14'b11100111111000;     //63pi/512
   cos[63]  =  14'b00111011010001;     //63pi/512
   sin[64]  =  14'b11100111100001;     //64pi/512
   cos[64]  =  14'b00111011001000;     //64pi/512
   sin[65]  =  14'b11100111001001;     //65pi/512
   cos[65]  =  14'b00111010111110;     //65pi/512
   sin[66]  =  14'b11100110110010;     //66pi/512
   cos[66]  =  14'b00111010110100;     //66pi/512
   sin[67]  =  14'b11100110011011;     //67pi/512
   cos[67]  =  14'b00111010101010;     //67pi/512
   sin[68]  =  14'b11100110000100;     //68pi/512
   cos[68]  =  14'b00111010100000;     //68pi/512
   sin[69]  =  14'b11100101101101;     //69pi/512
   cos[69]  =  14'b00111010010110;     //69pi/512
   sin[70]  =  14'b11100101010110;     //70pi/512
   cos[70]  =  14'b00111010001011;     //70pi/512
   sin[71]  =  14'b11100100111111;     //71pi/512
   cos[71]  =  14'b00111010000001;     //71pi/512
   sin[72]  =  14'b11100100101001;     //72pi/512
   cos[72]  =  14'b00111001110110;     //72pi/512
   sin[73]  =  14'b11100100010010;     //73pi/512
   cos[73]  =  14'b00111001101011;     //73pi/512
   sin[74]  =  14'b11100011111011;     //74pi/512
   cos[74]  =  14'b00111001100000;     //74pi/512
   sin[75]  =  14'b11100011100101;     //75pi/512
   cos[75]  =  14'b00111001010101;     //75pi/512
   sin[76]  =  14'b11100011001110;     //76pi/512
   cos[76]  =  14'b00111001001010;     //76pi/512
   sin[77]  =  14'b11100010111000;     //77pi/512
   cos[77]  =  14'b00111000111111;     //77pi/512
   sin[78]  =  14'b11100010100010;     //78pi/512
   cos[78]  =  14'b00111000110011;     //78pi/512
   sin[79]  =  14'b11100010001011;     //79pi/512
   cos[79]  =  14'b00111000101000;     //79pi/512
   sin[80]  =  14'b11100001110101;     //80pi/512
   cos[80]  =  14'b00111000011100;     //80pi/512
   sin[81]  =  14'b11100001011111;     //81pi/512
   cos[81]  =  14'b00111000010000;     //81pi/512
   sin[82]  =  14'b11100001001001;     //82pi/512
   cos[82]  =  14'b00111000000100;     //82pi/512
   sin[83]  =  14'b11100000110011;     //83pi/512
   cos[83]  =  14'b00110111111000;     //83pi/512
   sin[84]  =  14'b11100000011101;     //84pi/512
   cos[84]  =  14'b00110111101011;     //84pi/512
   sin[85]  =  14'b11100000000111;     //85pi/512
   cos[85]  =  14'b00110111011111;     //85pi/512
   sin[86]  =  14'b11011111110010;     //86pi/512
   cos[86]  =  14'b00110111010010;     //86pi/512
   sin[87]  =  14'b11011111011100;     //87pi/512
   cos[87]  =  14'b00110111000110;     //87pi/512
   sin[88]  =  14'b11011111000110;     //88pi/512
   cos[88]  =  14'b00110110111001;     //88pi/512
   sin[89]  =  14'b11011110110001;     //89pi/512
   cos[89]  =  14'b00110110101100;     //89pi/512
   sin[90]  =  14'b11011110011011;     //90pi/512
   cos[90]  =  14'b00110110011111;     //90pi/512
   sin[91]  =  14'b11011110000110;     //91pi/512
   cos[91]  =  14'b00110110010001;     //91pi/512
   sin[92]  =  14'b11011101110001;     //92pi/512
   cos[92]  =  14'b00110110000100;     //92pi/512
   sin[93]  =  14'b11011101011011;     //93pi/512
   cos[93]  =  14'b00110101110111;     //93pi/512
   sin[94]  =  14'b11011101000110;     //94pi/512
   cos[94]  =  14'b00110101101001;     //94pi/512
   sin[95]  =  14'b11011100110001;     //95pi/512
   cos[95]  =  14'b00110101011011;     //95pi/512
   sin[96]  =  14'b11011100011100;     //96pi/512
   cos[96]  =  14'b00110101001101;     //96pi/512
   sin[97]  =  14'b11011100001000;     //97pi/512
   cos[97]  =  14'b00110100111111;     //97pi/512
   sin[98]  =  14'b11011011110011;     //98pi/512
   cos[98]  =  14'b00110100110001;     //98pi/512
   sin[99]  =  14'b11011011011110;     //99pi/512
   cos[99]  =  14'b00110100100011;     //99pi/512
   sin[100]  =  14'b11011011001001;     //100pi/512
   cos[100]  =  14'b00110100010100;     //100pi/512
   sin[101]  =  14'b11011010110101;     //101pi/512
   cos[101]  =  14'b00110100000110;     //101pi/512
   sin[102]  =  14'b11011010100001;     //102pi/512
   cos[102]  =  14'b00110011110111;     //102pi/512
   sin[103]  =  14'b11011010001100;     //103pi/512
   cos[103]  =  14'b00110011101000;     //103pi/512
   sin[104]  =  14'b11011001111000;     //104pi/512
   cos[104]  =  14'b00110011011001;     //104pi/512
   sin[105]  =  14'b11011001100100;     //105pi/512
   cos[105]  =  14'b00110011001010;     //105pi/512
   sin[106]  =  14'b11011001010000;     //106pi/512
   cos[106]  =  14'b00110010111011;     //106pi/512
   sin[107]  =  14'b11011000111100;     //107pi/512
   cos[107]  =  14'b00110010101100;     //107pi/512
   sin[108]  =  14'b11011000101000;     //108pi/512
   cos[108]  =  14'b00110010011101;     //108pi/512
   sin[109]  =  14'b11011000010100;     //109pi/512
   cos[109]  =  14'b00110010001101;     //109pi/512
   sin[110]  =  14'b11011000000001;     //110pi/512
   cos[110]  =  14'b00110001111101;     //110pi/512
   sin[111]  =  14'b11010111101101;     //111pi/512
   cos[111]  =  14'b00110001101110;     //111pi/512
   sin[112]  =  14'b11010111011010;     //112pi/512
   cos[112]  =  14'b00110001011110;     //112pi/512
   sin[113]  =  14'b11010111000110;     //113pi/512
   cos[113]  =  14'b00110001001110;     //113pi/512
   sin[114]  =  14'b11010110110011;     //114pi/512
   cos[114]  =  14'b00110000111110;     //114pi/512
   sin[115]  =  14'b11010110100000;     //115pi/512
   cos[115]  =  14'b00110000101101;     //115pi/512
   sin[116]  =  14'b11010110001101;     //116pi/512
   cos[116]  =  14'b00110000011101;     //116pi/512
   sin[117]  =  14'b11010101111010;     //117pi/512
   cos[117]  =  14'b00110000001101;     //117pi/512
   sin[118]  =  14'b11010101100111;     //118pi/512
   cos[118]  =  14'b00101111111100;     //118pi/512
   sin[119]  =  14'b11010101010100;     //119pi/512
   cos[119]  =  14'b00101111101011;     //119pi/512
   sin[120]  =  14'b11010101000001;     //120pi/512
   cos[120]  =  14'b00101111011010;     //120pi/512
   sin[121]  =  14'b11010100101111;     //121pi/512
   cos[121]  =  14'b00101111001010;     //121pi/512
   sin[122]  =  14'b11010100011100;     //122pi/512
   cos[122]  =  14'b00101110111000;     //122pi/512
   sin[123]  =  14'b11010100001010;     //123pi/512
   cos[123]  =  14'b00101110100111;     //123pi/512
   sin[124]  =  14'b11010011111000;     //124pi/512
   cos[124]  =  14'b00101110010110;     //124pi/512
   sin[125]  =  14'b11010011100101;     //125pi/512
   cos[125]  =  14'b00101110000101;     //125pi/512
   sin[126]  =  14'b11010011010011;     //126pi/512
   cos[126]  =  14'b00101101110011;     //126pi/512
   sin[127]  =  14'b11010011000010;     //127pi/512
   cos[127]  =  14'b00101101100010;     //127pi/512
   sin[128]  =  14'b11010010110000;     //128pi/512
   cos[128]  =  14'b00101101010000;     //128pi/512
   sin[129]  =  14'b11010010011110;     //129pi/512
   cos[129]  =  14'b00101100111110;     //129pi/512
   sin[130]  =  14'b11010010001100;     //130pi/512
   cos[130]  =  14'b00101100101100;     //130pi/512
   sin[131]  =  14'b11010001111011;     //131pi/512
   cos[131]  =  14'b00101100011010;     //131pi/512
   sin[132]  =  14'b11010001101001;     //132pi/512
   cos[132]  =  14'b00101100001000;     //132pi/512
   sin[133]  =  14'b11010001011000;     //133pi/512
   cos[133]  =  14'b00101011110110;     //133pi/512
   sin[134]  =  14'b11010001000111;     //134pi/512
   cos[134]  =  14'b00101011100011;     //134pi/512
   sin[135]  =  14'b11010000110110;     //135pi/512
   cos[135]  =  14'b00101011010001;     //135pi/512
   sin[136]  =  14'b11010000100101;     //136pi/512
   cos[136]  =  14'b00101010111110;     //136pi/512
   sin[137]  =  14'b11010000010100;     //137pi/512
   cos[137]  =  14'b00101010101100;     //137pi/512
   sin[138]  =  14'b11010000000100;     //138pi/512
   cos[138]  =  14'b00101010011001;     //138pi/512
   sin[139]  =  14'b11001111110011;     //139pi/512
   cos[139]  =  14'b00101010000110;     //139pi/512
   sin[140]  =  14'b11001111100010;     //140pi/512
   cos[140]  =  14'b00101001110011;     //140pi/512
   sin[141]  =  14'b11001111010010;     //141pi/512
   cos[141]  =  14'b00101001100000;     //141pi/512
   sin[142]  =  14'b11001111000010;     //142pi/512
   cos[142]  =  14'b00101001001101;     //142pi/512
   sin[143]  =  14'b11001110110010;     //143pi/512
   cos[143]  =  14'b00101000111001;     //143pi/512
   sin[144]  =  14'b11001110100010;     //144pi/512
   cos[144]  =  14'b00101000100110;     //144pi/512
   sin[145]  =  14'b11001110010010;     //145pi/512
   cos[145]  =  14'b00101000010010;     //145pi/512
   sin[146]  =  14'b11001110000010;     //146pi/512
   cos[146]  =  14'b00100111111111;     //146pi/512
   sin[147]  =  14'b11001101110010;     //147pi/512
   cos[147]  =  14'b00100111101011;     //147pi/512
   sin[148]  =  14'b11001101100011;     //148pi/512
   cos[148]  =  14'b00100111010111;     //148pi/512
   sin[149]  =  14'b11001101010100;     //149pi/512
   cos[149]  =  14'b00100111000100;     //149pi/512
   sin[150]  =  14'b11001101000100;     //150pi/512
   cos[150]  =  14'b00100110110000;     //150pi/512
   sin[151]  =  14'b11001100110101;     //151pi/512
   cos[151]  =  14'b00100110011100;     //151pi/512
   sin[152]  =  14'b11001100100110;     //152pi/512
   cos[152]  =  14'b00100110000111;     //152pi/512
   sin[153]  =  14'b11001100010111;     //153pi/512
   cos[153]  =  14'b00100101110011;     //153pi/512
   sin[154]  =  14'b11001100001000;     //154pi/512
   cos[154]  =  14'b00100101011111;     //154pi/512
   sin[155]  =  14'b11001011111010;     //155pi/512
   cos[155]  =  14'b00100101001011;     //155pi/512
   sin[156]  =  14'b11001011101011;     //156pi/512
   cos[156]  =  14'b00100100110110;     //156pi/512
   sin[157]  =  14'b11001011011101;     //157pi/512
   cos[157]  =  14'b00100100100001;     //157pi/512
   sin[158]  =  14'b11001011001110;     //158pi/512
   cos[158]  =  14'b00100100001101;     //158pi/512
   sin[159]  =  14'b11001011000000;     //159pi/512
   cos[159]  =  14'b00100011111000;     //159pi/512
   sin[160]  =  14'b11001010110010;     //160pi/512
   cos[160]  =  14'b00100011100011;     //160pi/512
   sin[161]  =  14'b11001010100100;     //161pi/512
   cos[161]  =  14'b00100011001110;     //161pi/512
   sin[162]  =  14'b11001010010111;     //162pi/512
   cos[162]  =  14'b00100010111001;     //162pi/512
   sin[163]  =  14'b11001010001001;     //163pi/512
   cos[163]  =  14'b00100010100100;     //163pi/512
   sin[164]  =  14'b11001001111011;     //164pi/512
   cos[164]  =  14'b00100010001111;     //164pi/512
   sin[165]  =  14'b11001001101110;     //165pi/512
   cos[165]  =  14'b00100001111010;     //165pi/512
   sin[166]  =  14'b11001001100001;     //166pi/512
   cos[166]  =  14'b00100001100100;     //166pi/512
   sin[167]  =  14'b11001001010100;     //167pi/512
   cos[167]  =  14'b00100001001111;     //167pi/512
   sin[168]  =  14'b11001001000111;     //168pi/512
   cos[168]  =  14'b00100000111001;     //168pi/512
   sin[169]  =  14'b11001000111010;     //169pi/512
   cos[169]  =  14'b00100000100100;     //169pi/512
   sin[170]  =  14'b11001000101101;     //170pi/512
   cos[170]  =  14'b00100000001110;     //170pi/512
   sin[171]  =  14'b11001000100001;     //171pi/512
   cos[171]  =  14'b00011111111000;     //171pi/512
   sin[172]  =  14'b11001000010100;     //172pi/512
   cos[172]  =  14'b00011111100010;     //172pi/512
   sin[173]  =  14'b11001000001000;     //173pi/512
   cos[173]  =  14'b00011111001101;     //173pi/512
   sin[174]  =  14'b11000111111100;     //174pi/512
   cos[174]  =  14'b00011110110111;     //174pi/512
   sin[175]  =  14'b11000111110000;     //175pi/512
   cos[175]  =  14'b00011110100000;     //175pi/512
   sin[176]  =  14'b11000111100100;     //176pi/512
   cos[176]  =  14'b00011110001010;     //176pi/512
   sin[177]  =  14'b11000111011000;     //177pi/512
   cos[177]  =  14'b00011101110100;     //177pi/512
   sin[178]  =  14'b11000111001100;     //178pi/512
   cos[178]  =  14'b00011101011110;     //178pi/512
   sin[179]  =  14'b11000111000001;     //179pi/512
   cos[179]  =  14'b00011101001000;     //179pi/512
   sin[180]  =  14'b11000110110101;     //180pi/512
   cos[180]  =  14'b00011100110001;     //180pi/512
   sin[181]  =  14'b11000110101010;     //181pi/512
   cos[181]  =  14'b00011100011011;     //181pi/512
   sin[182]  =  14'b11000110011111;     //182pi/512
   cos[182]  =  14'b00011100000100;     //182pi/512
   sin[183]  =  14'b11000110010100;     //183pi/512
   cos[183]  =  14'b00011011101101;     //183pi/512
   sin[184]  =  14'b11000110001001;     //184pi/512
   cos[184]  =  14'b00011011010111;     //184pi/512
   sin[185]  =  14'b11000101111111;     //185pi/512
   cos[185]  =  14'b00011011000000;     //185pi/512
   sin[186]  =  14'b11000101110100;     //186pi/512
   cos[186]  =  14'b00011010101001;     //186pi/512
   sin[187]  =  14'b11000101101010;     //187pi/512
   cos[187]  =  14'b00011010010010;     //187pi/512
   sin[188]  =  14'b11000101011111;     //188pi/512
   cos[188]  =  14'b00011001111011;     //188pi/512
   sin[189]  =  14'b11000101010101;     //189pi/512
   cos[189]  =  14'b00011001100100;     //189pi/512
   sin[190]  =  14'b11000101001011;     //190pi/512
   cos[190]  =  14'b00011001001101;     //190pi/512
   sin[191]  =  14'b11000101000001;     //191pi/512
   cos[191]  =  14'b00011000110110;     //191pi/512
   sin[192]  =  14'b11000100111000;     //192pi/512
   cos[192]  =  14'b00011000011111;     //192pi/512
   sin[193]  =  14'b11000100101110;     //193pi/512
   cos[193]  =  14'b00011000001000;     //193pi/512
   sin[194]  =  14'b11000100100101;     //194pi/512
   cos[194]  =  14'b00010111110000;     //194pi/512
   sin[195]  =  14'b11000100011100;     //195pi/512
   cos[195]  =  14'b00010111011001;     //195pi/512
   sin[196]  =  14'b11000100010010;     //196pi/512
   cos[196]  =  14'b00010111000010;     //196pi/512
   sin[197]  =  14'b11000100001001;     //197pi/512
   cos[197]  =  14'b00010110101010;     //197pi/512
   sin[198]  =  14'b11000100000001;     //198pi/512
   cos[198]  =  14'b00010110010011;     //198pi/512
   sin[199]  =  14'b11000011111000;     //199pi/512
   cos[199]  =  14'b00010101111011;     //199pi/512
   sin[200]  =  14'b11000011101111;     //200pi/512
   cos[200]  =  14'b00010101100011;     //200pi/512
   sin[201]  =  14'b11000011100111;     //201pi/512
   cos[201]  =  14'b00010101001100;     //201pi/512
   sin[202]  =  14'b11000011011111;     //202pi/512
   cos[202]  =  14'b00010100110100;     //202pi/512
   sin[203]  =  14'b11000011010111;     //203pi/512
   cos[203]  =  14'b00010100011100;     //203pi/512
   sin[204]  =  14'b11000011001111;     //204pi/512
   cos[204]  =  14'b00010100000100;     //204pi/512
   sin[205]  =  14'b11000011000111;     //205pi/512
   cos[205]  =  14'b00010011101100;     //205pi/512
   sin[206]  =  14'b11000010111111;     //206pi/512
   cos[206]  =  14'b00010011010101;     //206pi/512
   sin[207]  =  14'b11000010111000;     //207pi/512
   cos[207]  =  14'b00010010111101;     //207pi/512
   sin[208]  =  14'b11000010110000;     //208pi/512
   cos[208]  =  14'b00010010100101;     //208pi/512
   sin[209]  =  14'b11000010101001;     //209pi/512
   cos[209]  =  14'b00010010001100;     //209pi/512
   sin[210]  =  14'b11000010100010;     //210pi/512
   cos[210]  =  14'b00010001110100;     //210pi/512
   sin[211]  =  14'b11000010011011;     //211pi/512
   cos[211]  =  14'b00010001011100;     //211pi/512
   sin[212]  =  14'b11000010010100;     //212pi/512
   cos[212]  =  14'b00010001000100;     //212pi/512
   sin[213]  =  14'b11000010001110;     //213pi/512
   cos[213]  =  14'b00010000101100;     //213pi/512
   sin[214]  =  14'b11000010000111;     //214pi/512
   cos[214]  =  14'b00010000010011;     //214pi/512
   sin[215]  =  14'b11000010000001;     //215pi/512
   cos[215]  =  14'b00001111111011;     //215pi/512
   sin[216]  =  14'b11000001111011;     //216pi/512
   cos[216]  =  14'b00001111100011;     //216pi/512
   sin[217]  =  14'b11000001110101;     //217pi/512
   cos[217]  =  14'b00001111001010;     //217pi/512
   sin[218]  =  14'b11000001101111;     //218pi/512
   cos[218]  =  14'b00001110110010;     //218pi/512
   sin[219]  =  14'b11000001101001;     //219pi/512
   cos[219]  =  14'b00001110011001;     //219pi/512
   sin[220]  =  14'b11000001100100;     //220pi/512
   cos[220]  =  14'b00001110000001;     //220pi/512
   sin[221]  =  14'b11000001011110;     //221pi/512
   cos[221]  =  14'b00001101101000;     //221pi/512
   sin[222]  =  14'b11000001011001;     //222pi/512
   cos[222]  =  14'b00001101010000;     //222pi/512
   sin[223]  =  14'b11000001010100;     //223pi/512
   cos[223]  =  14'b00001100110111;     //223pi/512
   sin[224]  =  14'b11000001001111;     //224pi/512
   cos[224]  =  14'b00001100011111;     //224pi/512
   sin[225]  =  14'b11000001001010;     //225pi/512
   cos[225]  =  14'b00001100000110;     //225pi/512
   sin[226]  =  14'b11000001000101;     //226pi/512
   cos[226]  =  14'b00001011101101;     //226pi/512
   sin[227]  =  14'b11000001000001;     //227pi/512
   cos[227]  =  14'b00001011010101;     //227pi/512
   sin[228]  =  14'b11000000111100;     //228pi/512
   cos[228]  =  14'b00001010111100;     //228pi/512
   sin[229]  =  14'b11000000111000;     //229pi/512
   cos[229]  =  14'b00001010100011;     //229pi/512
   sin[230]  =  14'b11000000110100;     //230pi/512
   cos[230]  =  14'b00001010001010;     //230pi/512
   sin[231]  =  14'b11000000110000;     //231pi/512
   cos[231]  =  14'b00001001110001;     //231pi/512
   sin[232]  =  14'b11000000101100;     //232pi/512
   cos[232]  =  14'b00001001011001;     //232pi/512
   sin[233]  =  14'b11000000101001;     //233pi/512
   cos[233]  =  14'b00001001000000;     //233pi/512
   sin[234]  =  14'b11000000100101;     //234pi/512
   cos[234]  =  14'b00001000100111;     //234pi/512
   sin[235]  =  14'b11000000100010;     //235pi/512
   cos[235]  =  14'b00001000001110;     //235pi/512
   sin[236]  =  14'b11000000011111;     //236pi/512
   cos[236]  =  14'b00000111110101;     //236pi/512
   sin[237]  =  14'b11000000011100;     //237pi/512
   cos[237]  =  14'b00000111011100;     //237pi/512
   sin[238]  =  14'b11000000011001;     //238pi/512
   cos[238]  =  14'b00000111000011;     //238pi/512
   sin[239]  =  14'b11000000010110;     //239pi/512
   cos[239]  =  14'b00000110101010;     //239pi/512
   sin[240]  =  14'b11000000010100;     //240pi/512
   cos[240]  =  14'b00000110010001;     //240pi/512
   sin[241]  =  14'b11000000010001;     //241pi/512
   cos[241]  =  14'b00000101111000;     //241pi/512
   sin[242]  =  14'b11000000001111;     //242pi/512
   cos[242]  =  14'b00000101011111;     //242pi/512
   sin[243]  =  14'b11000000001101;     //243pi/512
   cos[243]  =  14'b00000101000110;     //243pi/512
   sin[244]  =  14'b11000000001011;     //244pi/512
   cos[244]  =  14'b00000100101101;     //244pi/512
   sin[245]  =  14'b11000000001001;     //245pi/512
   cos[245]  =  14'b00000100010100;     //245pi/512
   sin[246]  =  14'b11000000001000;     //246pi/512
   cos[246]  =  14'b00000011111011;     //246pi/512
   sin[247]  =  14'b11000000000110;     //247pi/512
   cos[247]  =  14'b00000011100010;     //247pi/512
   sin[248]  =  14'b11000000000101;     //248pi/512
   cos[248]  =  14'b00000011001000;     //248pi/512
   sin[249]  =  14'b11000000000100;     //249pi/512
   cos[249]  =  14'b00000010101111;     //249pi/512
   sin[250]  =  14'b11000000000011;     //250pi/512
   cos[250]  =  14'b00000010010110;     //250pi/512
   sin[251]  =  14'b11000000000010;     //251pi/512
   cos[251]  =  14'b00000001111101;     //251pi/512
   sin[252]  =  14'b11000000000001;     //252pi/512
   cos[252]  =  14'b00000001100100;     //252pi/512
   sin[253]  =  14'b11000000000001;     //253pi/512
   cos[253]  =  14'b00000001001011;     //253pi/512
   sin[254]  =  14'b11000000000000;     //254pi/512
   cos[254]  =  14'b00000000110010;     //254pi/512
   sin[255]  =  14'b11000000000000;     //255pi/512
   cos[255]  =  14'b00000000011001;     //255pi/512
   sin[256]  =  14'b11000000000000;     //256pi/512
   cos[256]  =  14'b00000000000000;     //256pi/512
   sin[257]  =  14'b11000000000000;     //257pi/512
   cos[257]  =  14'b11111111100111;     //257pi/512
   sin[258]  =  14'b11000000000000;     //258pi/512
   cos[258]  =  14'b11111111001110;     //258pi/512
   sin[259]  =  14'b11000000000001;     //259pi/512
   cos[259]  =  14'b11111110110101;     //259pi/512
   sin[260]  =  14'b11000000000001;     //260pi/512
   cos[260]  =  14'b11111110011011;     //260pi/512
   sin[261]  =  14'b11000000000010;     //261pi/512
   cos[261]  =  14'b11111110000010;     //261pi/512
   sin[262]  =  14'b11000000000011;     //262pi/512
   cos[262]  =  14'b11111101101001;     //262pi/512
   sin[263]  =  14'b11000000000100;     //263pi/512
   cos[263]  =  14'b11111101010000;     //263pi/512
   sin[264]  =  14'b11000000000101;     //264pi/512
   cos[264]  =  14'b11111100110111;     //264pi/512
   sin[265]  =  14'b11000000000110;     //265pi/512
   cos[265]  =  14'b11111100011110;     //265pi/512
   sin[266]  =  14'b11000000001000;     //266pi/512
   cos[266]  =  14'b11111100000101;     //266pi/512
   sin[267]  =  14'b11000000001001;     //267pi/512
   cos[267]  =  14'b11111011101100;     //267pi/512
   sin[268]  =  14'b11000000001011;     //268pi/512
   cos[268]  =  14'b11111011010011;     //268pi/512
   sin[269]  =  14'b11000000001101;     //269pi/512
   cos[269]  =  14'b11111010111010;     //269pi/512
   sin[270]  =  14'b11000000001111;     //270pi/512
   cos[270]  =  14'b11111010100001;     //270pi/512
   sin[271]  =  14'b11000000010001;     //271pi/512
   cos[271]  =  14'b11111010001000;     //271pi/512
   sin[272]  =  14'b11000000010100;     //272pi/512
   cos[272]  =  14'b11111001101111;     //272pi/512
   sin[273]  =  14'b11000000010110;     //273pi/512
   cos[273]  =  14'b11111001010110;     //273pi/512
   sin[274]  =  14'b11000000011001;     //274pi/512
   cos[274]  =  14'b11111000111101;     //274pi/512
   sin[275]  =  14'b11000000011100;     //275pi/512
   cos[275]  =  14'b11111000100100;     //275pi/512
   sin[276]  =  14'b11000000011111;     //276pi/512
   cos[276]  =  14'b11111000001011;     //276pi/512
   sin[277]  =  14'b11000000100010;     //277pi/512
   cos[277]  =  14'b11110111110010;     //277pi/512
   sin[278]  =  14'b11000000100101;     //278pi/512
   cos[278]  =  14'b11110111011001;     //278pi/512
   sin[279]  =  14'b11000000101001;     //279pi/512
   cos[279]  =  14'b11110111000000;     //279pi/512
   sin[280]  =  14'b11000000101100;     //280pi/512
   cos[280]  =  14'b11110110100111;     //280pi/512
   sin[281]  =  14'b11000000110000;     //281pi/512
   cos[281]  =  14'b11110110001110;     //281pi/512
   sin[282]  =  14'b11000000110100;     //282pi/512
   cos[282]  =  14'b11110101110101;     //282pi/512
   sin[283]  =  14'b11000000111000;     //283pi/512
   cos[283]  =  14'b11110101011101;     //283pi/512
   sin[284]  =  14'b11000000111100;     //284pi/512
   cos[284]  =  14'b11110101000100;     //284pi/512
   sin[285]  =  14'b11000001000001;     //285pi/512
   cos[285]  =  14'b11110100101011;     //285pi/512
   sin[286]  =  14'b11000001000101;     //286pi/512
   cos[286]  =  14'b11110100010010;     //286pi/512
   sin[287]  =  14'b11000001001010;     //287pi/512
   cos[287]  =  14'b11110011111010;     //287pi/512
   sin[288]  =  14'b11000001001111;     //288pi/512
   cos[288]  =  14'b11110011100001;     //288pi/512
   sin[289]  =  14'b11000001010100;     //289pi/512
   cos[289]  =  14'b11110011001000;     //289pi/512
   sin[290]  =  14'b11000001011001;     //290pi/512
   cos[290]  =  14'b11110010110000;     //290pi/512
   sin[291]  =  14'b11000001011110;     //291pi/512
   cos[291]  =  14'b11110010010111;     //291pi/512
   sin[292]  =  14'b11000001100100;     //292pi/512
   cos[292]  =  14'b11110001111111;     //292pi/512
   sin[293]  =  14'b11000001101001;     //293pi/512
   cos[293]  =  14'b11110001100110;     //293pi/512
   sin[294]  =  14'b11000001101111;     //294pi/512
   cos[294]  =  14'b11110001001110;     //294pi/512
   sin[295]  =  14'b11000001110101;     //295pi/512
   cos[295]  =  14'b11110000110101;     //295pi/512
   sin[296]  =  14'b11000001111011;     //296pi/512
   cos[296]  =  14'b11110000011101;     //296pi/512
   sin[297]  =  14'b11000010000001;     //297pi/512
   cos[297]  =  14'b11110000000100;     //297pi/512
   sin[298]  =  14'b11000010000111;     //298pi/512
   cos[298]  =  14'b11101111101100;     //298pi/512
   sin[299]  =  14'b11000010001110;     //299pi/512
   cos[299]  =  14'b11101111010100;     //299pi/512
   sin[300]  =  14'b11000010010100;     //300pi/512
   cos[300]  =  14'b11101110111100;     //300pi/512
   sin[301]  =  14'b11000010011011;     //301pi/512
   cos[301]  =  14'b11101110100011;     //301pi/512
   sin[302]  =  14'b11000010100010;     //302pi/512
   cos[302]  =  14'b11101110001011;     //302pi/512
   sin[303]  =  14'b11000010101001;     //303pi/512
   cos[303]  =  14'b11101101110011;     //303pi/512
   sin[304]  =  14'b11000010110000;     //304pi/512
   cos[304]  =  14'b11101101011011;     //304pi/512
   sin[305]  =  14'b11000010111000;     //305pi/512
   cos[305]  =  14'b11101101000011;     //305pi/512
   sin[306]  =  14'b11000010111111;     //306pi/512
   cos[306]  =  14'b11101100101011;     //306pi/512
   sin[307]  =  14'b11000011000111;     //307pi/512
   cos[307]  =  14'b11101100010011;     //307pi/512
   sin[308]  =  14'b11000011001111;     //308pi/512
   cos[308]  =  14'b11101011111011;     //308pi/512
   sin[309]  =  14'b11000011010111;     //309pi/512
   cos[309]  =  14'b11101011100011;     //309pi/512
   sin[310]  =  14'b11000011011111;     //310pi/512
   cos[310]  =  14'b11101011001100;     //310pi/512
   sin[311]  =  14'b11000011100111;     //311pi/512
   cos[311]  =  14'b11101010110100;     //311pi/512
   sin[312]  =  14'b11000011101111;     //312pi/512
   cos[312]  =  14'b11101010011100;     //312pi/512
   sin[313]  =  14'b11000011111000;     //313pi/512
   cos[313]  =  14'b11101010000100;     //313pi/512
   sin[314]  =  14'b11000100000001;     //314pi/512
   cos[314]  =  14'b11101001101101;     //314pi/512
   sin[315]  =  14'b11000100001001;     //315pi/512
   cos[315]  =  14'b11101001010101;     //315pi/512
   sin[316]  =  14'b11000100010010;     //316pi/512
   cos[316]  =  14'b11101000111110;     //316pi/512
   sin[317]  =  14'b11000100011100;     //317pi/512
   cos[317]  =  14'b11101000100110;     //317pi/512
   sin[318]  =  14'b11000100100101;     //318pi/512
   cos[318]  =  14'b11101000001111;     //318pi/512
   sin[319]  =  14'b11000100101110;     //319pi/512
   cos[319]  =  14'b11100111111000;     //319pi/512
   sin[320]  =  14'b11000100111000;     //320pi/512
   cos[320]  =  14'b11100111100001;     //320pi/512
   sin[321]  =  14'b11000101000001;     //321pi/512
   cos[321]  =  14'b11100111001001;     //321pi/512
   sin[322]  =  14'b11000101001011;     //322pi/512
   cos[322]  =  14'b11100110110010;     //322pi/512
   sin[323]  =  14'b11000101010101;     //323pi/512
   cos[323]  =  14'b11100110011011;     //323pi/512
   sin[324]  =  14'b11000101011111;     //324pi/512
   cos[324]  =  14'b11100110000100;     //324pi/512
   sin[325]  =  14'b11000101101010;     //325pi/512
   cos[325]  =  14'b11100101101101;     //325pi/512
   sin[326]  =  14'b11000101110100;     //326pi/512
   cos[326]  =  14'b11100101010110;     //326pi/512
   sin[327]  =  14'b11000101111111;     //327pi/512
   cos[327]  =  14'b11100100111111;     //327pi/512
   sin[328]  =  14'b11000110001001;     //328pi/512
   cos[328]  =  14'b11100100101001;     //328pi/512
   sin[329]  =  14'b11000110010100;     //329pi/512
   cos[329]  =  14'b11100100010010;     //329pi/512
   sin[330]  =  14'b11000110011111;     //330pi/512
   cos[330]  =  14'b11100011111011;     //330pi/512
   sin[331]  =  14'b11000110101010;     //331pi/512
   cos[331]  =  14'b11100011100101;     //331pi/512
   sin[332]  =  14'b11000110110101;     //332pi/512
   cos[332]  =  14'b11100011001110;     //332pi/512
   sin[333]  =  14'b11000111000001;     //333pi/512
   cos[333]  =  14'b11100010111000;     //333pi/512
   sin[334]  =  14'b11000111001100;     //334pi/512
   cos[334]  =  14'b11100010100010;     //334pi/512
   sin[335]  =  14'b11000111011000;     //335pi/512
   cos[335]  =  14'b11100010001011;     //335pi/512
   sin[336]  =  14'b11000111100100;     //336pi/512
   cos[336]  =  14'b11100001110101;     //336pi/512
   sin[337]  =  14'b11000111110000;     //337pi/512
   cos[337]  =  14'b11100001011111;     //337pi/512
   sin[338]  =  14'b11000111111100;     //338pi/512
   cos[338]  =  14'b11100001001001;     //338pi/512
   sin[339]  =  14'b11001000001000;     //339pi/512
   cos[339]  =  14'b11100000110011;     //339pi/512
   sin[340]  =  14'b11001000010100;     //340pi/512
   cos[340]  =  14'b11100000011101;     //340pi/512
   sin[341]  =  14'b11001000100001;     //341pi/512
   cos[341]  =  14'b11100000000111;     //341pi/512
   sin[342]  =  14'b11001000101101;     //342pi/512
   cos[342]  =  14'b11011111110010;     //342pi/512
   sin[343]  =  14'b11001000111010;     //343pi/512
   cos[343]  =  14'b11011111011100;     //343pi/512
   sin[344]  =  14'b11001001000111;     //344pi/512
   cos[344]  =  14'b11011111000110;     //344pi/512
   sin[345]  =  14'b11001001010100;     //345pi/512
   cos[345]  =  14'b11011110110001;     //345pi/512
   sin[346]  =  14'b11001001100001;     //346pi/512
   cos[346]  =  14'b11011110011011;     //346pi/512
   sin[347]  =  14'b11001001101110;     //347pi/512
   cos[347]  =  14'b11011110000110;     //347pi/512
   sin[348]  =  14'b11001001111011;     //348pi/512
   cos[348]  =  14'b11011101110001;     //348pi/512
   sin[349]  =  14'b11001010001001;     //349pi/512
   cos[349]  =  14'b11011101011011;     //349pi/512
   sin[350]  =  14'b11001010010111;     //350pi/512
   cos[350]  =  14'b11011101000110;     //350pi/512
   sin[351]  =  14'b11001010100100;     //351pi/512
   cos[351]  =  14'b11011100110001;     //351pi/512
   sin[352]  =  14'b11001010110010;     //352pi/512
   cos[352]  =  14'b11011100011100;     //352pi/512
   sin[353]  =  14'b11001011000000;     //353pi/512
   cos[353]  =  14'b11011100001000;     //353pi/512
   sin[354]  =  14'b11001011001110;     //354pi/512
   cos[354]  =  14'b11011011110011;     //354pi/512
   sin[355]  =  14'b11001011011101;     //355pi/512
   cos[355]  =  14'b11011011011110;     //355pi/512
   sin[356]  =  14'b11001011101011;     //356pi/512
   cos[356]  =  14'b11011011001001;     //356pi/512
   sin[357]  =  14'b11001011111010;     //357pi/512
   cos[357]  =  14'b11011010110101;     //357pi/512
   sin[358]  =  14'b11001100001000;     //358pi/512
   cos[358]  =  14'b11011010100001;     //358pi/512
   sin[359]  =  14'b11001100010111;     //359pi/512
   cos[359]  =  14'b11011010001100;     //359pi/512
   sin[360]  =  14'b11001100100110;     //360pi/512
   cos[360]  =  14'b11011001111000;     //360pi/512
   sin[361]  =  14'b11001100110101;     //361pi/512
   cos[361]  =  14'b11011001100100;     //361pi/512
   sin[362]  =  14'b11001101000100;     //362pi/512
   cos[362]  =  14'b11011001010000;     //362pi/512
   sin[363]  =  14'b11001101010100;     //363pi/512
   cos[363]  =  14'b11011000111100;     //363pi/512
   sin[364]  =  14'b11001101100011;     //364pi/512
   cos[364]  =  14'b11011000101000;     //364pi/512
   sin[365]  =  14'b11001101110010;     //365pi/512
   cos[365]  =  14'b11011000010100;     //365pi/512
   sin[366]  =  14'b11001110000010;     //366pi/512
   cos[366]  =  14'b11011000000001;     //366pi/512
   sin[367]  =  14'b11001110010010;     //367pi/512
   cos[367]  =  14'b11010111101101;     //367pi/512
   sin[368]  =  14'b11001110100010;     //368pi/512
   cos[368]  =  14'b11010111011010;     //368pi/512
   sin[369]  =  14'b11001110110010;     //369pi/512
   cos[369]  =  14'b11010111000110;     //369pi/512
   sin[370]  =  14'b11001111000010;     //370pi/512
   cos[370]  =  14'b11010110110011;     //370pi/512
   sin[371]  =  14'b11001111010010;     //371pi/512
   cos[371]  =  14'b11010110100000;     //371pi/512
   sin[372]  =  14'b11001111100010;     //372pi/512
   cos[372]  =  14'b11010110001101;     //372pi/512
   sin[373]  =  14'b11001111110011;     //373pi/512
   cos[373]  =  14'b11010101111010;     //373pi/512
   sin[374]  =  14'b11010000000100;     //374pi/512
   cos[374]  =  14'b11010101100111;     //374pi/512
   sin[375]  =  14'b11010000010100;     //375pi/512
   cos[375]  =  14'b11010101010100;     //375pi/512
   sin[376]  =  14'b11010000100101;     //376pi/512
   cos[376]  =  14'b11010101000001;     //376pi/512
   sin[377]  =  14'b11010000110110;     //377pi/512
   cos[377]  =  14'b11010100101111;     //377pi/512
   sin[378]  =  14'b11010001000111;     //378pi/512
   cos[378]  =  14'b11010100011100;     //378pi/512
   sin[379]  =  14'b11010001011000;     //379pi/512
   cos[379]  =  14'b11010100001010;     //379pi/512
   sin[380]  =  14'b11010001101001;     //380pi/512
   cos[380]  =  14'b11010011111000;     //380pi/512
   sin[381]  =  14'b11010001111011;     //381pi/512
   cos[381]  =  14'b11010011100101;     //381pi/512
   sin[382]  =  14'b11010010001100;     //382pi/512
   cos[382]  =  14'b11010011010011;     //382pi/512
   sin[383]  =  14'b11010010011110;     //383pi/512
   cos[383]  =  14'b11010011000010;     //383pi/512
   sin[384]  =  14'b11010010110000;     //384pi/512
   cos[384]  =  14'b11010010110000;     //384pi/512
   sin[385]  =  14'b11010011000010;     //385pi/512
   cos[385]  =  14'b11010010011110;     //385pi/512
   sin[386]  =  14'b11010011010011;     //386pi/512
   cos[386]  =  14'b11010010001100;     //386pi/512
   sin[387]  =  14'b11010011100101;     //387pi/512
   cos[387]  =  14'b11010001111011;     //387pi/512
   sin[388]  =  14'b11010011111000;     //388pi/512
   cos[388]  =  14'b11010001101001;     //388pi/512
   sin[389]  =  14'b11010100001010;     //389pi/512
   cos[389]  =  14'b11010001011000;     //389pi/512
   sin[390]  =  14'b11010100011100;     //390pi/512
   cos[390]  =  14'b11010001000111;     //390pi/512
   sin[391]  =  14'b11010100101111;     //391pi/512
   cos[391]  =  14'b11010000110110;     //391pi/512
   sin[392]  =  14'b11010101000001;     //392pi/512
   cos[392]  =  14'b11010000100101;     //392pi/512
   sin[393]  =  14'b11010101010100;     //393pi/512
   cos[393]  =  14'b11010000010100;     //393pi/512
   sin[394]  =  14'b11010101100111;     //394pi/512
   cos[394]  =  14'b11010000000100;     //394pi/512
   sin[395]  =  14'b11010101111010;     //395pi/512
   cos[395]  =  14'b11001111110011;     //395pi/512
   sin[396]  =  14'b11010110001101;     //396pi/512
   cos[396]  =  14'b11001111100010;     //396pi/512
   sin[397]  =  14'b11010110100000;     //397pi/512
   cos[397]  =  14'b11001111010010;     //397pi/512
   sin[398]  =  14'b11010110110011;     //398pi/512
   cos[398]  =  14'b11001111000010;     //398pi/512
   sin[399]  =  14'b11010111000110;     //399pi/512
   cos[399]  =  14'b11001110110010;     //399pi/512
   sin[400]  =  14'b11010111011010;     //400pi/512
   cos[400]  =  14'b11001110100010;     //400pi/512
   sin[401]  =  14'b11010111101101;     //401pi/512
   cos[401]  =  14'b11001110010010;     //401pi/512
   sin[402]  =  14'b11011000000001;     //402pi/512
   cos[402]  =  14'b11001110000010;     //402pi/512
   sin[403]  =  14'b11011000010100;     //403pi/512
   cos[403]  =  14'b11001101110010;     //403pi/512
   sin[404]  =  14'b11011000101000;     //404pi/512
   cos[404]  =  14'b11001101100011;     //404pi/512
   sin[405]  =  14'b11011000111100;     //405pi/512
   cos[405]  =  14'b11001101010100;     //405pi/512
   sin[406]  =  14'b11011001010000;     //406pi/512
   cos[406]  =  14'b11001101000100;     //406pi/512
   sin[407]  =  14'b11011001100100;     //407pi/512
   cos[407]  =  14'b11001100110101;     //407pi/512
   sin[408]  =  14'b11011001111000;     //408pi/512
   cos[408]  =  14'b11001100100110;     //408pi/512
   sin[409]  =  14'b11011010001100;     //409pi/512
   cos[409]  =  14'b11001100010111;     //409pi/512
   sin[410]  =  14'b11011010100001;     //410pi/512
   cos[410]  =  14'b11001100001000;     //410pi/512
   sin[411]  =  14'b11011010110101;     //411pi/512
   cos[411]  =  14'b11001011111010;     //411pi/512
   sin[412]  =  14'b11011011001001;     //412pi/512
   cos[412]  =  14'b11001011101011;     //412pi/512
   sin[413]  =  14'b11011011011110;     //413pi/512
   cos[413]  =  14'b11001011011101;     //413pi/512
   sin[414]  =  14'b11011011110011;     //414pi/512
   cos[414]  =  14'b11001011001110;     //414pi/512
   sin[415]  =  14'b11011100001000;     //415pi/512
   cos[415]  =  14'b11001011000000;     //415pi/512
   sin[416]  =  14'b11011100011100;     //416pi/512
   cos[416]  =  14'b11001010110010;     //416pi/512
   sin[417]  =  14'b11011100110001;     //417pi/512
   cos[417]  =  14'b11001010100100;     //417pi/512
   sin[418]  =  14'b11011101000110;     //418pi/512
   cos[418]  =  14'b11001010010111;     //418pi/512
   sin[419]  =  14'b11011101011011;     //419pi/512
   cos[419]  =  14'b11001010001001;     //419pi/512
   sin[420]  =  14'b11011101110001;     //420pi/512
   cos[420]  =  14'b11001001111011;     //420pi/512
   sin[421]  =  14'b11011110000110;     //421pi/512
   cos[421]  =  14'b11001001101110;     //421pi/512
   sin[422]  =  14'b11011110011011;     //422pi/512
   cos[422]  =  14'b11001001100001;     //422pi/512
   sin[423]  =  14'b11011110110001;     //423pi/512
   cos[423]  =  14'b11001001010100;     //423pi/512
   sin[424]  =  14'b11011111000110;     //424pi/512
   cos[424]  =  14'b11001001000111;     //424pi/512
   sin[425]  =  14'b11011111011100;     //425pi/512
   cos[425]  =  14'b11001000111010;     //425pi/512
   sin[426]  =  14'b11011111110010;     //426pi/512
   cos[426]  =  14'b11001000101101;     //426pi/512
   sin[427]  =  14'b11100000000111;     //427pi/512
   cos[427]  =  14'b11001000100001;     //427pi/512
   sin[428]  =  14'b11100000011101;     //428pi/512
   cos[428]  =  14'b11001000010100;     //428pi/512
   sin[429]  =  14'b11100000110011;     //429pi/512
   cos[429]  =  14'b11001000001000;     //429pi/512
   sin[430]  =  14'b11100001001001;     //430pi/512
   cos[430]  =  14'b11000111111100;     //430pi/512
   sin[431]  =  14'b11100001011111;     //431pi/512
   cos[431]  =  14'b11000111110000;     //431pi/512
   sin[432]  =  14'b11100001110101;     //432pi/512
   cos[432]  =  14'b11000111100100;     //432pi/512
   sin[433]  =  14'b11100010001011;     //433pi/512
   cos[433]  =  14'b11000111011000;     //433pi/512
   sin[434]  =  14'b11100010100010;     //434pi/512
   cos[434]  =  14'b11000111001100;     //434pi/512
   sin[435]  =  14'b11100010111000;     //435pi/512
   cos[435]  =  14'b11000111000001;     //435pi/512
   sin[436]  =  14'b11100011001110;     //436pi/512
   cos[436]  =  14'b11000110110101;     //436pi/512
   sin[437]  =  14'b11100011100101;     //437pi/512
   cos[437]  =  14'b11000110101010;     //437pi/512
   sin[438]  =  14'b11100011111011;     //438pi/512
   cos[438]  =  14'b11000110011111;     //438pi/512
   sin[439]  =  14'b11100100010010;     //439pi/512
   cos[439]  =  14'b11000110010100;     //439pi/512
   sin[440]  =  14'b11100100101001;     //440pi/512
   cos[440]  =  14'b11000110001001;     //440pi/512
   sin[441]  =  14'b11100100111111;     //441pi/512
   cos[441]  =  14'b11000101111111;     //441pi/512
   sin[442]  =  14'b11100101010110;     //442pi/512
   cos[442]  =  14'b11000101110100;     //442pi/512
   sin[443]  =  14'b11100101101101;     //443pi/512
   cos[443]  =  14'b11000101101010;     //443pi/512
   sin[444]  =  14'b11100110000100;     //444pi/512
   cos[444]  =  14'b11000101011111;     //444pi/512
   sin[445]  =  14'b11100110011011;     //445pi/512
   cos[445]  =  14'b11000101010101;     //445pi/512
   sin[446]  =  14'b11100110110010;     //446pi/512
   cos[446]  =  14'b11000101001011;     //446pi/512
   sin[447]  =  14'b11100111001001;     //447pi/512
   cos[447]  =  14'b11000101000001;     //447pi/512
   sin[448]  =  14'b11100111100001;     //448pi/512
   cos[448]  =  14'b11000100111000;     //448pi/512
   sin[449]  =  14'b11100111111000;     //449pi/512
   cos[449]  =  14'b11000100101110;     //449pi/512
   sin[450]  =  14'b11101000001111;     //450pi/512
   cos[450]  =  14'b11000100100101;     //450pi/512
   sin[451]  =  14'b11101000100110;     //451pi/512
   cos[451]  =  14'b11000100011100;     //451pi/512
   sin[452]  =  14'b11101000111110;     //452pi/512
   cos[452]  =  14'b11000100010010;     //452pi/512
   sin[453]  =  14'b11101001010101;     //453pi/512
   cos[453]  =  14'b11000100001001;     //453pi/512
   sin[454]  =  14'b11101001101101;     //454pi/512
   cos[454]  =  14'b11000100000001;     //454pi/512
   sin[455]  =  14'b11101010000100;     //455pi/512
   cos[455]  =  14'b11000011111000;     //455pi/512
   sin[456]  =  14'b11101010011100;     //456pi/512
   cos[456]  =  14'b11000011101111;     //456pi/512
   sin[457]  =  14'b11101010110100;     //457pi/512
   cos[457]  =  14'b11000011100111;     //457pi/512
   sin[458]  =  14'b11101011001100;     //458pi/512
   cos[458]  =  14'b11000011011111;     //458pi/512
   sin[459]  =  14'b11101011100011;     //459pi/512
   cos[459]  =  14'b11000011010111;     //459pi/512
   sin[460]  =  14'b11101011111011;     //460pi/512
   cos[460]  =  14'b11000011001111;     //460pi/512
   sin[461]  =  14'b11101100010011;     //461pi/512
   cos[461]  =  14'b11000011000111;     //461pi/512
   sin[462]  =  14'b11101100101011;     //462pi/512
   cos[462]  =  14'b11000010111111;     //462pi/512
   sin[463]  =  14'b11101101000011;     //463pi/512
   cos[463]  =  14'b11000010111000;     //463pi/512
   sin[464]  =  14'b11101101011011;     //464pi/512
   cos[464]  =  14'b11000010110000;     //464pi/512
   sin[465]  =  14'b11101101110011;     //465pi/512
   cos[465]  =  14'b11000010101001;     //465pi/512
   sin[466]  =  14'b11101110001011;     //466pi/512
   cos[466]  =  14'b11000010100010;     //466pi/512
   sin[467]  =  14'b11101110100011;     //467pi/512
   cos[467]  =  14'b11000010011011;     //467pi/512
   sin[468]  =  14'b11101110111100;     //468pi/512
   cos[468]  =  14'b11000010010100;     //468pi/512
   sin[469]  =  14'b11101111010100;     //469pi/512
   cos[469]  =  14'b11000010001110;     //469pi/512
   sin[470]  =  14'b11101111101100;     //470pi/512
   cos[470]  =  14'b11000010000111;     //470pi/512
   sin[471]  =  14'b11110000000100;     //471pi/512
   cos[471]  =  14'b11000010000001;     //471pi/512
   sin[472]  =  14'b11110000011101;     //472pi/512
   cos[472]  =  14'b11000001111011;     //472pi/512
   sin[473]  =  14'b11110000110101;     //473pi/512
   cos[473]  =  14'b11000001110101;     //473pi/512
   sin[474]  =  14'b11110001001110;     //474pi/512
   cos[474]  =  14'b11000001101111;     //474pi/512
   sin[475]  =  14'b11110001100110;     //475pi/512
   cos[475]  =  14'b11000001101001;     //475pi/512
   sin[476]  =  14'b11110001111111;     //476pi/512
   cos[476]  =  14'b11000001100100;     //476pi/512
   sin[477]  =  14'b11110010010111;     //477pi/512
   cos[477]  =  14'b11000001011110;     //477pi/512
   sin[478]  =  14'b11110010110000;     //478pi/512
   cos[478]  =  14'b11000001011001;     //478pi/512
   sin[479]  =  14'b11110011001000;     //479pi/512
   cos[479]  =  14'b11000001010100;     //479pi/512
   sin[480]  =  14'b11110011100001;     //480pi/512
   cos[480]  =  14'b11000001001111;     //480pi/512
   sin[481]  =  14'b11110011111010;     //481pi/512
   cos[481]  =  14'b11000001001010;     //481pi/512
   sin[482]  =  14'b11110100010010;     //482pi/512
   cos[482]  =  14'b11000001000101;     //482pi/512
   sin[483]  =  14'b11110100101011;     //483pi/512
   cos[483]  =  14'b11000001000001;     //483pi/512
   sin[484]  =  14'b11110101000100;     //484pi/512
   cos[484]  =  14'b11000000111100;     //484pi/512
   sin[485]  =  14'b11110101011101;     //485pi/512
   cos[485]  =  14'b11000000111000;     //485pi/512
   sin[486]  =  14'b11110101110101;     //486pi/512
   cos[486]  =  14'b11000000110100;     //486pi/512
   sin[487]  =  14'b11110110001110;     //487pi/512
   cos[487]  =  14'b11000000110000;     //487pi/512
   sin[488]  =  14'b11110110100111;     //488pi/512
   cos[488]  =  14'b11000000101100;     //488pi/512
   sin[489]  =  14'b11110111000000;     //489pi/512
   cos[489]  =  14'b11000000101001;     //489pi/512
   sin[490]  =  14'b11110111011001;     //490pi/512
   cos[490]  =  14'b11000000100101;     //490pi/512
   sin[491]  =  14'b11110111110010;     //491pi/512
   cos[491]  =  14'b11000000100010;     //491pi/512
   sin[492]  =  14'b11111000001011;     //492pi/512
   cos[492]  =  14'b11000000011111;     //492pi/512
   sin[493]  =  14'b11111000100100;     //493pi/512
   cos[493]  =  14'b11000000011100;     //493pi/512
   sin[494]  =  14'b11111000111101;     //494pi/512
   cos[494]  =  14'b11000000011001;     //494pi/512
   sin[495]  =  14'b11111001010110;     //495pi/512
   cos[495]  =  14'b11000000010110;     //495pi/512
   sin[496]  =  14'b11111001101111;     //496pi/512
   cos[496]  =  14'b11000000010100;     //496pi/512
   sin[497]  =  14'b11111010001000;     //497pi/512
   cos[497]  =  14'b11000000010001;     //497pi/512
   sin[498]  =  14'b11111010100001;     //498pi/512
   cos[498]  =  14'b11000000001111;     //498pi/512
   sin[499]  =  14'b11111010111010;     //499pi/512
   cos[499]  =  14'b11000000001101;     //499pi/512
   sin[500]  =  14'b11111011010011;     //500pi/512
   cos[500]  =  14'b11000000001011;     //500pi/512
   sin[501]  =  14'b11111011101100;     //501pi/512
   cos[501]  =  14'b11000000001001;     //501pi/512
   sin[502]  =  14'b11111100000101;     //502pi/512
   cos[502]  =  14'b11000000001000;     //502pi/512
   sin[503]  =  14'b11111100011110;     //503pi/512
   cos[503]  =  14'b11000000000110;     //503pi/512
   sin[504]  =  14'b11111100110111;     //504pi/512
   cos[504]  =  14'b11000000000101;     //504pi/512
   sin[505]  =  14'b11111101010000;     //505pi/512
   cos[505]  =  14'b11000000000100;     //505pi/512
   sin[506]  =  14'b11111101101001;     //506pi/512
   cos[506]  =  14'b11000000000011;     //506pi/512
   sin[507]  =  14'b11111110000010;     //507pi/512
   cos[507]  =  14'b11000000000010;     //507pi/512
   sin[508]  =  14'b11111110011011;     //508pi/512
   cos[508]  =  14'b11000000000001;     //508pi/512
   sin[509]  =  14'b11111110110101;     //509pi/512
   cos[509]  =  14'b11000000000001;     //509pi/512
   sin[510]  =  14'b11111111001110;     //510pi/512
   cos[510]  =  14'b11000000000000;     //510pi/512
   sin[511]  =  14'b11111111100111;     //511pi/512
   cos[511]  =  14'b11000000000000;     //511pi/512

   sin[512]  =  14'b00000000000000;     //0pi/512
   cos[512]  =  14'b01000000000000;     //0pi/512
   sin[513]  =  14'b11111111101100;     //1pi/512
   cos[513]  =  14'b00111111111111;     //1pi/512
   sin[514]  =  14'b11111111011000;     //2pi/512
   cos[514]  =  14'b00111111111111;     //2pi/512
   sin[515]  =  14'b11111111000100;     //3pi/512
   cos[515]  =  14'b00111111111111;     //3pi/512
   sin[516]  =  14'b11111110110000;     //4pi/512
   cos[516]  =  14'b00111111111111;     //4pi/512
   sin[517]  =  14'b11111110011011;     //5pi/512
   cos[517]  =  14'b00111111111110;     //5pi/512
   sin[518]  =  14'b11111110000111;     //6pi/512
   cos[518]  =  14'b00111111111110;     //6pi/512
   sin[519]  =  14'b11111101110011;     //7pi/512
   cos[519]  =  14'b00111111111101;     //7pi/512
   sin[520]  =  14'b11111101011111;     //8pi/512
   cos[520]  =  14'b00111111111100;     //8pi/512
   sin[521]  =  14'b11111101001011;     //9pi/512
   cos[521]  =  14'b00111111111100;     //9pi/512
   sin[522]  =  14'b11111100110111;     //10pi/512
   cos[522]  =  14'b00111111111011;     //10pi/512
   sin[523]  =  14'b11111100100011;     //11pi/512
   cos[523]  =  14'b00111111111010;     //11pi/512
   sin[524]  =  14'b11111100001111;     //12pi/512
   cos[524]  =  14'b00111111111000;     //12pi/512
   sin[525]  =  14'b11111011111011;     //13pi/512
   cos[525]  =  14'b00111111110111;     //13pi/512
   sin[526]  =  14'b11111011100111;     //14pi/512
   cos[526]  =  14'b00111111110110;     //14pi/512
   sin[527]  =  14'b11111011010011;     //15pi/512
   cos[527]  =  14'b00111111110100;     //15pi/512
   sin[528]  =  14'b11111010111111;     //16pi/512
   cos[528]  =  14'b00111111110011;     //16pi/512
   sin[529]  =  14'b11111010101011;     //17pi/512
   cos[529]  =  14'b00111111110001;     //17pi/512
   sin[530]  =  14'b11111010010111;     //18pi/512
   cos[530]  =  14'b00111111110000;     //18pi/512
   sin[531]  =  14'b11111010000011;     //19pi/512
   cos[531]  =  14'b00111111101110;     //19pi/512
   sin[532]  =  14'b11111001101111;     //20pi/512
   cos[532]  =  14'b00111111101100;     //20pi/512
   sin[533]  =  14'b11111001011011;     //21pi/512
   cos[533]  =  14'b00111111101010;     //21pi/512
   sin[534]  =  14'b11111001000111;     //22pi/512
   cos[534]  =  14'b00111111101000;     //22pi/512
   sin[535]  =  14'b11111000110011;     //23pi/512
   cos[535]  =  14'b00111111100101;     //23pi/512
   sin[536]  =  14'b11111000011111;     //24pi/512
   cos[536]  =  14'b00111111100011;     //24pi/512
   sin[537]  =  14'b11111000001011;     //25pi/512
   cos[537]  =  14'b00111111100001;     //25pi/512
   sin[538]  =  14'b11110111110111;     //26pi/512
   cos[538]  =  14'b00111111011110;     //26pi/512
   sin[539]  =  14'b11110111100011;     //27pi/512
   cos[539]  =  14'b00111111011100;     //27pi/512
   sin[540]  =  14'b11110111001111;     //28pi/512
   cos[540]  =  14'b00111111011001;     //28pi/512
   sin[541]  =  14'b11110110111011;     //29pi/512
   cos[541]  =  14'b00111111010110;     //29pi/512
   sin[542]  =  14'b11110110100111;     //30pi/512
   cos[542]  =  14'b00111111010011;     //30pi/512
   sin[543]  =  14'b11110110010011;     //31pi/512
   cos[543]  =  14'b00111111010000;     //31pi/512
   sin[544]  =  14'b11110101111111;     //32pi/512
   cos[544]  =  14'b00111111001101;     //32pi/512
   sin[545]  =  14'b11110101101011;     //33pi/512
   cos[545]  =  14'b00111111001010;     //33pi/512
   sin[546]  =  14'b11110101011000;     //34pi/512
   cos[546]  =  14'b00111111000111;     //34pi/512
   sin[547]  =  14'b11110101000100;     //35pi/512
   cos[547]  =  14'b00111111000011;     //35pi/512
   sin[548]  =  14'b11110100110000;     //36pi/512
   cos[548]  =  14'b00111111000000;     //36pi/512
   sin[549]  =  14'b11110100011100;     //37pi/512
   cos[549]  =  14'b00111110111100;     //37pi/512
   sin[550]  =  14'b11110100001000;     //38pi/512
   cos[550]  =  14'b00111110111000;     //38pi/512
   sin[551]  =  14'b11110011110101;     //39pi/512
   cos[551]  =  14'b00111110110101;     //39pi/512
   sin[552]  =  14'b11110011100001;     //40pi/512
   cos[552]  =  14'b00111110110001;     //40pi/512
   sin[553]  =  14'b11110011001101;     //41pi/512
   cos[553]  =  14'b00111110101101;     //41pi/512
   sin[554]  =  14'b11110010111010;     //42pi/512
   cos[554]  =  14'b00111110101001;     //42pi/512
   sin[555]  =  14'b11110010100110;     //43pi/512
   cos[555]  =  14'b00111110100101;     //43pi/512
   sin[556]  =  14'b11110010010010;     //44pi/512
   cos[556]  =  14'b00111110100000;     //44pi/512
   sin[557]  =  14'b11110001111111;     //45pi/512
   cos[557]  =  14'b00111110011100;     //45pi/512
   sin[558]  =  14'b11110001101011;     //46pi/512
   cos[558]  =  14'b00111110011000;     //46pi/512
   sin[559]  =  14'b11110001010111;     //47pi/512
   cos[559]  =  14'b00111110010011;     //47pi/512
   sin[560]  =  14'b11110001000100;     //48pi/512
   cos[560]  =  14'b00111110001110;     //48pi/512
   sin[561]  =  14'b11110000110000;     //49pi/512
   cos[561]  =  14'b00111110001010;     //49pi/512
   sin[562]  =  14'b11110000011101;     //50pi/512
   cos[562]  =  14'b00111110000101;     //50pi/512
   sin[563]  =  14'b11110000001001;     //51pi/512
   cos[563]  =  14'b00111110000000;     //51pi/512
   sin[564]  =  14'b11101111110110;     //52pi/512
   cos[564]  =  14'b00111101111011;     //52pi/512
   sin[565]  =  14'b11101111100010;     //53pi/512
   cos[565]  =  14'b00111101110110;     //53pi/512
   sin[566]  =  14'b11101111001111;     //54pi/512
   cos[566]  =  14'b00111101110000;     //54pi/512
   sin[567]  =  14'b11101110111100;     //55pi/512
   cos[567]  =  14'b00111101101011;     //55pi/512
   sin[568]  =  14'b11101110101000;     //56pi/512
   cos[568]  =  14'b00111101100110;     //56pi/512
   sin[569]  =  14'b11101110010101;     //57pi/512
   cos[569]  =  14'b00111101100000;     //57pi/512
   sin[570]  =  14'b11101110000010;     //58pi/512
   cos[570]  =  14'b00111101011011;     //58pi/512
   sin[571]  =  14'b11101101101110;     //59pi/512
   cos[571]  =  14'b00111101010101;     //59pi/512
   sin[572]  =  14'b11101101011011;     //60pi/512
   cos[572]  =  14'b00111101001111;     //60pi/512
   sin[573]  =  14'b11101101001000;     //61pi/512
   cos[573]  =  14'b00111101001001;     //61pi/512
   sin[574]  =  14'b11101100110101;     //62pi/512
   cos[574]  =  14'b00111101000011;     //62pi/512
   sin[575]  =  14'b11101100100001;     //63pi/512
   cos[575]  =  14'b00111100111101;     //63pi/512
   sin[576]  =  14'b11101100001110;     //64pi/512
   cos[576]  =  14'b00111100110111;     //64pi/512
   sin[577]  =  14'b11101011111011;     //65pi/512
   cos[577]  =  14'b00111100110001;     //65pi/512
   sin[578]  =  14'b11101011101000;     //66pi/512
   cos[578]  =  14'b00111100101010;     //66pi/512
   sin[579]  =  14'b11101011010101;     //67pi/512
   cos[579]  =  14'b00111100100100;     //67pi/512
   sin[580]  =  14'b11101011000010;     //68pi/512
   cos[580]  =  14'b00111100011101;     //68pi/512
   sin[581]  =  14'b11101010101111;     //69pi/512
   cos[581]  =  14'b00111100010111;     //69pi/512
   sin[582]  =  14'b11101010011100;     //70pi/512
   cos[582]  =  14'b00111100010000;     //70pi/512
   sin[583]  =  14'b11101010001001;     //71pi/512
   cos[583]  =  14'b00111100001001;     //71pi/512
   sin[584]  =  14'b11101001110110;     //72pi/512
   cos[584]  =  14'b00111100000010;     //72pi/512
   sin[585]  =  14'b11101001100011;     //73pi/512
   cos[585]  =  14'b00111011111011;     //73pi/512
   sin[586]  =  14'b11101001010001;     //74pi/512
   cos[586]  =  14'b00111011110100;     //74pi/512
   sin[587]  =  14'b11101000111110;     //75pi/512
   cos[587]  =  14'b00111011101101;     //75pi/512
   sin[588]  =  14'b11101000101011;     //76pi/512
   cos[588]  =  14'b00111011100110;     //76pi/512
   sin[589]  =  14'b11101000011000;     //77pi/512
   cos[589]  =  14'b00111011011110;     //77pi/512
   sin[590]  =  14'b11101000000110;     //78pi/512
   cos[590]  =  14'b00111011010111;     //78pi/512
   sin[591]  =  14'b11100111110011;     //79pi/512
   cos[591]  =  14'b00111011001111;     //79pi/512
   sin[592]  =  14'b11100111100001;     //80pi/512
   cos[592]  =  14'b00111011001000;     //80pi/512
   sin[593]  =  14'b11100111001110;     //81pi/512
   cos[593]  =  14'b00111011000000;     //81pi/512
   sin[594]  =  14'b11100110111011;     //82pi/512
   cos[594]  =  14'b00111010111000;     //82pi/512
   sin[595]  =  14'b11100110101001;     //83pi/512
   cos[595]  =  14'b00111010110000;     //83pi/512
   sin[596]  =  14'b11100110010111;     //84pi/512
   cos[596]  =  14'b00111010101000;     //84pi/512
   sin[597]  =  14'b11100110000100;     //85pi/512
   cos[597]  =  14'b00111010100000;     //85pi/512
   sin[598]  =  14'b11100101110010;     //86pi/512
   cos[598]  =  14'b00111010011000;     //86pi/512
   sin[599]  =  14'b11100101011111;     //87pi/512
   cos[599]  =  14'b00111010010000;     //87pi/512
   sin[600]  =  14'b11100101001101;     //88pi/512
   cos[600]  =  14'b00111010000111;     //88pi/512
   sin[601]  =  14'b11100100111011;     //89pi/512
   cos[601]  =  14'b00111001111111;     //89pi/512
   sin[602]  =  14'b11100100101001;     //90pi/512
   cos[602]  =  14'b00111001110110;     //90pi/512
   sin[603]  =  14'b11100100010111;     //91pi/512
   cos[603]  =  14'b00111001101110;     //91pi/512
   sin[604]  =  14'b11100100000100;     //92pi/512
   cos[604]  =  14'b00111001100101;     //92pi/512
   sin[605]  =  14'b11100011110010;     //93pi/512
   cos[605]  =  14'b00111001011100;     //93pi/512
   sin[606]  =  14'b11100011100000;     //94pi/512
   cos[606]  =  14'b00111001010011;     //94pi/512
   sin[607]  =  14'b11100011001110;     //95pi/512
   cos[607]  =  14'b00111001001010;     //95pi/512
   sin[608]  =  14'b11100010111100;     //96pi/512
   cos[608]  =  14'b00111001000001;     //96pi/512
   sin[609]  =  14'b11100010101011;     //97pi/512
   cos[609]  =  14'b00111000111000;     //97pi/512
   sin[610]  =  14'b11100010011001;     //98pi/512
   cos[610]  =  14'b00111000101111;     //98pi/512
   sin[611]  =  14'b11100010000111;     //99pi/512
   cos[611]  =  14'b00111000100101;     //99pi/512
   sin[612]  =  14'b11100001110101;     //100pi/512
   cos[612]  =  14'b00111000011100;     //100pi/512
   sin[613]  =  14'b11100001100011;     //101pi/512
   cos[613]  =  14'b00111000010010;     //101pi/512
   sin[614]  =  14'b11100001010010;     //102pi/512
   cos[614]  =  14'b00111000001001;     //102pi/512
   sin[615]  =  14'b11100001000000;     //103pi/512
   cos[615]  =  14'b00110111111111;     //103pi/512
   sin[616]  =  14'b11100000101111;     //104pi/512
   cos[616]  =  14'b00110111110101;     //104pi/512
   sin[617]  =  14'b11100000011101;     //105pi/512
   cos[617]  =  14'b00110111101011;     //105pi/512
   sin[618]  =  14'b11100000001100;     //106pi/512
   cos[618]  =  14'b00110111100001;     //106pi/512
   sin[619]  =  14'b11011111111010;     //107pi/512
   cos[619]  =  14'b00110111010111;     //107pi/512
   sin[620]  =  14'b11011111101001;     //108pi/512
   cos[620]  =  14'b00110111001101;     //108pi/512
   sin[621]  =  14'b11011111011000;     //109pi/512
   cos[621]  =  14'b00110111000011;     //109pi/512
   sin[622]  =  14'b11011111000110;     //110pi/512
   cos[622]  =  14'b00110110111001;     //110pi/512
   sin[623]  =  14'b11011110110101;     //111pi/512
   cos[623]  =  14'b00110110101110;     //111pi/512
   sin[624]  =  14'b11011110100100;     //112pi/512
   cos[624]  =  14'b00110110100100;     //112pi/512
   sin[625]  =  14'b11011110010011;     //113pi/512
   cos[625]  =  14'b00110110011001;     //113pi/512
   sin[626]  =  14'b11011110000010;     //114pi/512
   cos[626]  =  14'b00110110001111;     //114pi/512
   sin[627]  =  14'b11011101110001;     //115pi/512
   cos[627]  =  14'b00110110000100;     //115pi/512
   sin[628]  =  14'b11011101100000;     //116pi/512
   cos[628]  =  14'b00110101111001;     //116pi/512
   sin[629]  =  14'b11011101001111;     //117pi/512
   cos[629]  =  14'b00110101101110;     //117pi/512
   sin[630]  =  14'b11011100111110;     //118pi/512
   cos[630]  =  14'b00110101100011;     //118pi/512
   sin[631]  =  14'b11011100101101;     //119pi/512
   cos[631]  =  14'b00110101011000;     //119pi/512
   sin[632]  =  14'b11011100011100;     //120pi/512
   cos[632]  =  14'b00110101001101;     //120pi/512
   sin[633]  =  14'b11011100001100;     //121pi/512
   cos[633]  =  14'b00110101000010;     //121pi/512
   sin[634]  =  14'b11011011111011;     //122pi/512
   cos[634]  =  14'b00110100110111;     //122pi/512
   sin[635]  =  14'b11011011101010;     //123pi/512
   cos[635]  =  14'b00110100101011;     //123pi/512
   sin[636]  =  14'b11011011011010;     //124pi/512
   cos[636]  =  14'b00110100100000;     //124pi/512
   sin[637]  =  14'b11011011001001;     //125pi/512
   cos[637]  =  14'b00110100010100;     //125pi/512
   sin[638]  =  14'b11011010111001;     //126pi/512
   cos[638]  =  14'b00110100001001;     //126pi/512
   sin[639]  =  14'b11011010101001;     //127pi/512
   cos[639]  =  14'b00110011111101;     //127pi/512
   sin[640]  =  14'b11011010011000;     //128pi/512
   cos[640]  =  14'b00110011110001;     //128pi/512
   sin[641]  =  14'b11011010001000;     //129pi/512
   cos[641]  =  14'b00110011100101;     //129pi/512
   sin[642]  =  14'b11011001111000;     //130pi/512
   cos[642]  =  14'b00110011011001;     //130pi/512
   sin[643]  =  14'b11011001101000;     //131pi/512
   cos[643]  =  14'b00110011001101;     //131pi/512
   sin[644]  =  14'b11011001011000;     //132pi/512
   cos[644]  =  14'b00110011000001;     //132pi/512
   sin[645]  =  14'b11011001001000;     //133pi/512
   cos[645]  =  14'b00110010110101;     //133pi/512
   sin[646]  =  14'b11011000111000;     //134pi/512
   cos[646]  =  14'b00110010101001;     //134pi/512
   sin[647]  =  14'b11011000101000;     //135pi/512
   cos[647]  =  14'b00110010011101;     //135pi/512
   sin[648]  =  14'b11011000011000;     //136pi/512
   cos[648]  =  14'b00110010010000;     //136pi/512
   sin[649]  =  14'b11011000001000;     //137pi/512
   cos[649]  =  14'b00110010000100;     //137pi/512
   sin[650]  =  14'b11010111111001;     //138pi/512
   cos[650]  =  14'b00110001110111;     //138pi/512
   sin[651]  =  14'b11010111101001;     //139pi/512
   cos[651]  =  14'b00110001101010;     //139pi/512
   sin[652]  =  14'b11010111011010;     //140pi/512
   cos[652]  =  14'b00110001011110;     //140pi/512
   sin[653]  =  14'b11010111001010;     //141pi/512
   cos[653]  =  14'b00110001010001;     //141pi/512
   sin[654]  =  14'b11010110111011;     //142pi/512
   cos[654]  =  14'b00110001000100;     //142pi/512
   sin[655]  =  14'b11010110101011;     //143pi/512
   cos[655]  =  14'b00110000110111;     //143pi/512
   sin[656]  =  14'b11010110011100;     //144pi/512
   cos[656]  =  14'b00110000101010;     //144pi/512
   sin[657]  =  14'b11010110001101;     //145pi/512
   cos[657]  =  14'b00110000011101;     //145pi/512
   sin[658]  =  14'b11010101111101;     //146pi/512
   cos[658]  =  14'b00110000010000;     //146pi/512
   sin[659]  =  14'b11010101101110;     //147pi/512
   cos[659]  =  14'b00110000000011;     //147pi/512
   sin[660]  =  14'b11010101011111;     //148pi/512
   cos[660]  =  14'b00101111110101;     //148pi/512
   sin[661]  =  14'b11010101010000;     //149pi/512
   cos[661]  =  14'b00101111101000;     //149pi/512
   sin[662]  =  14'b11010101000001;     //150pi/512
   cos[662]  =  14'b00101111011010;     //150pi/512
   sin[663]  =  14'b11010100110010;     //151pi/512
   cos[663]  =  14'b00101111001101;     //151pi/512
   sin[664]  =  14'b11010100100100;     //152pi/512
   cos[664]  =  14'b00101110111111;     //152pi/512
   sin[665]  =  14'b11010100010101;     //153pi/512
   cos[665]  =  14'b00101110110010;     //153pi/512
   sin[666]  =  14'b11010100000110;     //154pi/512
   cos[666]  =  14'b00101110100100;     //154pi/512
   sin[667]  =  14'b11010011111000;     //155pi/512
   cos[667]  =  14'b00101110010110;     //155pi/512
   sin[668]  =  14'b11010011101001;     //156pi/512
   cos[668]  =  14'b00101110001000;     //156pi/512
   sin[669]  =  14'b11010011011011;     //157pi/512
   cos[669]  =  14'b00101101111010;     //157pi/512
   sin[670]  =  14'b11010011001100;     //158pi/512
   cos[670]  =  14'b00101101101100;     //158pi/512
   sin[671]  =  14'b11010010111110;     //159pi/512
   cos[671]  =  14'b00101101011110;     //159pi/512
   sin[672]  =  14'b11010010110000;     //160pi/512
   cos[672]  =  14'b00101101010000;     //160pi/512
   sin[673]  =  14'b11010010100010;     //161pi/512
   cos[673]  =  14'b00101101000010;     //161pi/512
   sin[674]  =  14'b11010010010011;     //162pi/512
   cos[674]  =  14'b00101100110011;     //162pi/512
   sin[675]  =  14'b11010010000101;     //163pi/512
   cos[675]  =  14'b00101100100101;     //163pi/512
   sin[676]  =  14'b11010001110111;     //164pi/512
   cos[676]  =  14'b00101100010110;     //164pi/512
   sin[677]  =  14'b11010001101001;     //165pi/512
   cos[677]  =  14'b00101100001000;     //165pi/512
   sin[678]  =  14'b11010001011100;     //166pi/512
   cos[678]  =  14'b00101011111001;     //166pi/512
   sin[679]  =  14'b11010001001110;     //167pi/512
   cos[679]  =  14'b00101011101011;     //167pi/512
   sin[680]  =  14'b11010001000000;     //168pi/512
   cos[680]  =  14'b00101011011100;     //168pi/512
   sin[681]  =  14'b11010000110011;     //169pi/512
   cos[681]  =  14'b00101011001101;     //169pi/512
   sin[682]  =  14'b11010000100101;     //170pi/512
   cos[682]  =  14'b00101010111110;     //170pi/512
   sin[683]  =  14'b11010000011000;     //171pi/512
   cos[683]  =  14'b00101010101111;     //171pi/512
   sin[684]  =  14'b11010000001010;     //172pi/512
   cos[684]  =  14'b00101010100000;     //172pi/512
   sin[685]  =  14'b11001111111101;     //173pi/512
   cos[685]  =  14'b00101010010001;     //173pi/512
   sin[686]  =  14'b11001111110000;     //174pi/512
   cos[686]  =  14'b00101010000010;     //174pi/512
   sin[687]  =  14'b11001111100010;     //175pi/512
   cos[687]  =  14'b00101001110011;     //175pi/512
   sin[688]  =  14'b11001111010101;     //176pi/512
   cos[688]  =  14'b00101001100100;     //176pi/512
   sin[689]  =  14'b11001111001000;     //177pi/512
   cos[689]  =  14'b00101001010100;     //177pi/512
   sin[690]  =  14'b11001110111011;     //178pi/512
   cos[690]  =  14'b00101001000101;     //178pi/512
   sin[691]  =  14'b11001110101111;     //179pi/512
   cos[691]  =  14'b00101000110101;     //179pi/512
   sin[692]  =  14'b11001110100010;     //180pi/512
   cos[692]  =  14'b00101000100110;     //180pi/512
   sin[693]  =  14'b11001110010101;     //181pi/512
   cos[693]  =  14'b00101000010110;     //181pi/512
   sin[694]  =  14'b11001110001000;     //182pi/512
   cos[694]  =  14'b00101000000111;     //182pi/512
   sin[695]  =  14'b11001101111100;     //183pi/512
   cos[695]  =  14'b00100111110111;     //183pi/512
   sin[696]  =  14'b11001101101111;     //184pi/512
   cos[696]  =  14'b00100111100111;     //184pi/512
   sin[697]  =  14'b11001101100011;     //185pi/512
   cos[697]  =  14'b00100111010111;     //185pi/512
   sin[698]  =  14'b11001101010111;     //186pi/512
   cos[698]  =  14'b00100111001000;     //186pi/512
   sin[699]  =  14'b11001101001010;     //187pi/512
   cos[699]  =  14'b00100110111000;     //187pi/512
   sin[700]  =  14'b11001100111110;     //188pi/512
   cos[700]  =  14'b00100110101000;     //188pi/512
   sin[701]  =  14'b11001100110010;     //189pi/512
   cos[701]  =  14'b00100110011000;     //189pi/512
   sin[702]  =  14'b11001100100110;     //190pi/512
   cos[702]  =  14'b00100110000111;     //190pi/512
   sin[703]  =  14'b11001100011010;     //191pi/512
   cos[703]  =  14'b00100101110111;     //191pi/512
   sin[704]  =  14'b11001100001110;     //192pi/512
   cos[704]  =  14'b00100101100111;     //192pi/512
   sin[705]  =  14'b11001100000010;     //193pi/512
   cos[705]  =  14'b00100101010111;     //193pi/512
   sin[706]  =  14'b11001011110111;     //194pi/512
   cos[706]  =  14'b00100101000110;     //194pi/512
   sin[707]  =  14'b11001011101011;     //195pi/512
   cos[707]  =  14'b00100100110110;     //195pi/512
   sin[708]  =  14'b11001011100000;     //196pi/512
   cos[708]  =  14'b00100100100110;     //196pi/512
   sin[709]  =  14'b11001011010100;     //197pi/512
   cos[709]  =  14'b00100100010101;     //197pi/512
   sin[710]  =  14'b11001011001001;     //198pi/512
   cos[710]  =  14'b00100100000100;     //198pi/512
   sin[711]  =  14'b11001010111110;     //199pi/512
   cos[711]  =  14'b00100011110100;     //199pi/512
   sin[712]  =  14'b11001010110010;     //200pi/512
   cos[712]  =  14'b00100011100011;     //200pi/512
   sin[713]  =  14'b11001010100111;     //201pi/512
   cos[713]  =  14'b00100011010010;     //201pi/512
   sin[714]  =  14'b11001010011100;     //202pi/512
   cos[714]  =  14'b00100011000010;     //202pi/512
   sin[715]  =  14'b11001010010001;     //203pi/512
   cos[715]  =  14'b00100010110001;     //203pi/512
   sin[716]  =  14'b11001010000110;     //204pi/512
   cos[716]  =  14'b00100010100000;     //204pi/512
   sin[717]  =  14'b11001001111011;     //205pi/512
   cos[717]  =  14'b00100010001111;     //205pi/512
   sin[718]  =  14'b11001001110001;     //206pi/512
   cos[718]  =  14'b00100001111110;     //206pi/512
   sin[719]  =  14'b11001001100110;     //207pi/512
   cos[719]  =  14'b00100001101101;     //207pi/512
   sin[720]  =  14'b11001001011100;     //208pi/512
   cos[720]  =  14'b00100001011100;     //208pi/512
   sin[721]  =  14'b11001001010001;     //209pi/512
   cos[721]  =  14'b00100001001010;     //209pi/512
   sin[722]  =  14'b11001001000111;     //210pi/512
   cos[722]  =  14'b00100000111001;     //210pi/512
   sin[723]  =  14'b11001000111100;     //211pi/512
   cos[723]  =  14'b00100000101000;     //211pi/512
   sin[724]  =  14'b11001000110010;     //212pi/512
   cos[724]  =  14'b00100000010111;     //212pi/512
   sin[725]  =  14'b11001000101000;     //213pi/512
   cos[725]  =  14'b00100000000101;     //213pi/512
   sin[726]  =  14'b11001000011110;     //214pi/512
   cos[726]  =  14'b00011111110100;     //214pi/512
   sin[727]  =  14'b11001000010100;     //215pi/512
   cos[727]  =  14'b00011111100010;     //215pi/512
   sin[728]  =  14'b11001000001010;     //216pi/512
   cos[728]  =  14'b00011111010001;     //216pi/512
   sin[729]  =  14'b11001000000000;     //217pi/512
   cos[729]  =  14'b00011110111111;     //217pi/512
   sin[730]  =  14'b11000111110111;     //218pi/512
   cos[730]  =  14'b00011110101110;     //218pi/512
   sin[731]  =  14'b11000111101101;     //219pi/512
   cos[731]  =  14'b00011110011100;     //219pi/512
   sin[732]  =  14'b11000111100100;     //220pi/512
   cos[732]  =  14'b00011110001010;     //220pi/512
   sin[733]  =  14'b11000111011010;     //221pi/512
   cos[733]  =  14'b00011101111001;     //221pi/512
   sin[734]  =  14'b11000111010001;     //222pi/512
   cos[734]  =  14'b00011101100111;     //222pi/512
   sin[735]  =  14'b11000111001000;     //223pi/512
   cos[735]  =  14'b00011101010101;     //223pi/512
   sin[736]  =  14'b11000110111110;     //224pi/512
   cos[736]  =  14'b00011101000011;     //224pi/512
   sin[737]  =  14'b11000110110101;     //225pi/512
   cos[737]  =  14'b00011100110001;     //225pi/512
   sin[738]  =  14'b11000110101100;     //226pi/512
   cos[738]  =  14'b00011100011111;     //226pi/512
   sin[739]  =  14'b11000110100011;     //227pi/512
   cos[739]  =  14'b00011100001101;     //227pi/512
   sin[740]  =  14'b11000110011011;     //228pi/512
   cos[740]  =  14'b00011011111011;     //228pi/512
   sin[741]  =  14'b11000110010010;     //229pi/512
   cos[741]  =  14'b00011011101001;     //229pi/512
   sin[742]  =  14'b11000110001001;     //230pi/512
   cos[742]  =  14'b00011011010111;     //230pi/512
   sin[743]  =  14'b11000110000001;     //231pi/512
   cos[743]  =  14'b00011011000101;     //231pi/512
   sin[744]  =  14'b11000101111000;     //232pi/512
   cos[744]  =  14'b00011010110010;     //232pi/512
   sin[745]  =  14'b11000101110000;     //233pi/512
   cos[745]  =  14'b00011010100000;     //233pi/512
   sin[746]  =  14'b11000101101000;     //234pi/512
   cos[746]  =  14'b00011010001110;     //234pi/512
   sin[747]  =  14'b11000101011111;     //235pi/512
   cos[747]  =  14'b00011001111011;     //235pi/512
   sin[748]  =  14'b11000101010111;     //236pi/512
   cos[748]  =  14'b00011001101001;     //236pi/512
   sin[749]  =  14'b11000101001111;     //237pi/512
   cos[749]  =  14'b00011001010111;     //237pi/512
   sin[750]  =  14'b11000101000111;     //238pi/512
   cos[750]  =  14'b00011001000100;     //238pi/512
   sin[751]  =  14'b11000101000000;     //239pi/512
   cos[751]  =  14'b00011000110010;     //239pi/512
   sin[752]  =  14'b11000100111000;     //240pi/512
   cos[752]  =  14'b00011000011111;     //240pi/512
   sin[753]  =  14'b11000100110000;     //241pi/512
   cos[753]  =  14'b00011000001100;     //241pi/512
   sin[754]  =  14'b11000100101001;     //242pi/512
   cos[754]  =  14'b00010111111010;     //242pi/512
   sin[755]  =  14'b11000100100001;     //243pi/512
   cos[755]  =  14'b00010111100111;     //243pi/512
   sin[756]  =  14'b11000100011010;     //244pi/512
   cos[756]  =  14'b00010111010100;     //244pi/512
   sin[757]  =  14'b11000100010010;     //245pi/512
   cos[757]  =  14'b00010111000010;     //245pi/512
   sin[758]  =  14'b11000100001011;     //246pi/512
   cos[758]  =  14'b00010110101111;     //246pi/512
   sin[759]  =  14'b11000100000100;     //247pi/512
   cos[759]  =  14'b00010110011100;     //247pi/512
   sin[760]  =  14'b11000011111101;     //248pi/512
   cos[760]  =  14'b00010110001001;     //248pi/512
   sin[761]  =  14'b11000011110110;     //249pi/512
   cos[761]  =  14'b00010101110110;     //249pi/512
   sin[762]  =  14'b11000011101111;     //250pi/512
   cos[762]  =  14'b00010101100011;     //250pi/512
   sin[763]  =  14'b11000011101001;     //251pi/512
   cos[763]  =  14'b00010101010000;     //251pi/512
   sin[764]  =  14'b11000011100010;     //252pi/512
   cos[764]  =  14'b00010100111101;     //252pi/512
   sin[765]  =  14'b11000011011100;     //253pi/512
   cos[765]  =  14'b00010100101010;     //253pi/512
   sin[766]  =  14'b11000011010101;     //254pi/512
   cos[766]  =  14'b00010100010111;     //254pi/512
   sin[767]  =  14'b11000011001111;     //255pi/512
   cos[767]  =  14'b00010100000100;     //255pi/512
   sin[768]  =  14'b11000011001000;     //256pi/512
   cos[768]  =  14'b00010011110001;     //256pi/512
   sin[769]  =  14'b11000011000010;     //257pi/512
   cos[769]  =  14'b00010011011110;     //257pi/512
   sin[770]  =  14'b11000010111100;     //258pi/512
   cos[770]  =  14'b00010011001011;     //258pi/512
   sin[771]  =  14'b11000010110110;     //259pi/512
   cos[771]  =  14'b00010010111000;     //259pi/512
   sin[772]  =  14'b11000010110000;     //260pi/512
   cos[772]  =  14'b00010010100101;     //260pi/512
   sin[773]  =  14'b11000010101011;     //261pi/512
   cos[773]  =  14'b00010010010001;     //261pi/512
   sin[774]  =  14'b11000010100101;     //262pi/512
   cos[774]  =  14'b00010001111110;     //262pi/512
   sin[775]  =  14'b11000010011111;     //263pi/512
   cos[775]  =  14'b00010001101011;     //263pi/512
   sin[776]  =  14'b11000010011010;     //264pi/512
   cos[776]  =  14'b00010001010111;     //264pi/512
   sin[777]  =  14'b11000010010100;     //265pi/512
   cos[777]  =  14'b00010001000100;     //265pi/512
   sin[778]  =  14'b11000010001111;     //266pi/512
   cos[778]  =  14'b00010000110001;     //266pi/512
   sin[779]  =  14'b11000010001010;     //267pi/512
   cos[779]  =  14'b00010000011101;     //267pi/512
   sin[780]  =  14'b11000010000101;     //268pi/512
   cos[780]  =  14'b00010000001010;     //268pi/512
   sin[781]  =  14'b11000010000000;     //269pi/512
   cos[781]  =  14'b00001111110110;     //269pi/512
   sin[782]  =  14'b11000001111011;     //270pi/512
   cos[782]  =  14'b00001111100011;     //270pi/512
   sin[783]  =  14'b11000001110110;     //271pi/512
   cos[783]  =  14'b00001111001111;     //271pi/512
   sin[784]  =  14'b11000001110001;     //272pi/512
   cos[784]  =  14'b00001110111100;     //272pi/512
   sin[785]  =  14'b11000001101101;     //273pi/512
   cos[785]  =  14'b00001110101000;     //273pi/512
   sin[786]  =  14'b11000001101000;     //274pi/512
   cos[786]  =  14'b00001110010101;     //274pi/512
   sin[787]  =  14'b11000001100100;     //275pi/512
   cos[787]  =  14'b00001110000001;     //275pi/512
   sin[788]  =  14'b11000001011111;     //276pi/512
   cos[788]  =  14'b00001101101101;     //276pi/512
   sin[789]  =  14'b11000001011011;     //277pi/512
   cos[789]  =  14'b00001101011010;     //277pi/512
   sin[790]  =  14'b11000001010111;     //278pi/512
   cos[790]  =  14'b00001101000110;     //278pi/512
   sin[791]  =  14'b11000001010011;     //279pi/512
   cos[791]  =  14'b00001100110010;     //279pi/512
   sin[792]  =  14'b11000001001111;     //280pi/512
   cos[792]  =  14'b00001100011111;     //280pi/512
   sin[793]  =  14'b11000001001011;     //281pi/512
   cos[793]  =  14'b00001100001011;     //281pi/512
   sin[794]  =  14'b11000001000111;     //282pi/512
   cos[794]  =  14'b00001011110111;     //282pi/512
   sin[795]  =  14'b11000001000011;     //283pi/512
   cos[795]  =  14'b00001011100011;     //283pi/512
   sin[796]  =  14'b11000001000000;     //284pi/512
   cos[796]  =  14'b00001011010000;     //284pi/512
   sin[797]  =  14'b11000000111100;     //285pi/512
   cos[797]  =  14'b00001010111100;     //285pi/512
   sin[798]  =  14'b11000000111001;     //286pi/512
   cos[798]  =  14'b00001010101000;     //286pi/512
   sin[799]  =  14'b11000000110110;     //287pi/512
   cos[799]  =  14'b00001010010100;     //287pi/512
   sin[800]  =  14'b11000000110010;     //288pi/512
   cos[800]  =  14'b00001010000000;     //288pi/512
   sin[801]  =  14'b11000000101111;     //289pi/512
   cos[801]  =  14'b00001001101100;     //289pi/512
   sin[802]  =  14'b11000000101100;     //290pi/512
   cos[802]  =  14'b00001001011001;     //290pi/512
   sin[803]  =  14'b11000000101001;     //291pi/512
   cos[803]  =  14'b00001001000101;     //291pi/512
   sin[804]  =  14'b11000000100111;     //292pi/512
   cos[804]  =  14'b00001000110001;     //292pi/512
   sin[805]  =  14'b11000000100100;     //293pi/512
   cos[805]  =  14'b00001000011101;     //293pi/512
   sin[806]  =  14'b11000000100001;     //294pi/512
   cos[806]  =  14'b00001000001001;     //294pi/512
   sin[807]  =  14'b11000000011111;     //295pi/512
   cos[807]  =  14'b00000111110101;     //295pi/512
   sin[808]  =  14'b11000000011100;     //296pi/512
   cos[808]  =  14'b00000111100001;     //296pi/512
   sin[809]  =  14'b11000000011010;     //297pi/512
   cos[809]  =  14'b00000111001101;     //297pi/512
   sin[810]  =  14'b11000000011000;     //298pi/512
   cos[810]  =  14'b00000110111001;     //298pi/512
   sin[811]  =  14'b11000000010110;     //299pi/512
   cos[811]  =  14'b00000110100101;     //299pi/512
   sin[812]  =  14'b11000000010100;     //300pi/512
   cos[812]  =  14'b00000110010001;     //300pi/512
   sin[813]  =  14'b11000000010010;     //301pi/512
   cos[813]  =  14'b00000101111101;     //301pi/512
   sin[814]  =  14'b11000000010000;     //302pi/512
   cos[814]  =  14'b00000101101001;     //302pi/512
   sin[815]  =  14'b11000000001110;     //303pi/512
   cos[815]  =  14'b00000101010101;     //303pi/512
   sin[816]  =  14'b11000000001101;     //304pi/512
   cos[816]  =  14'b00000101000001;     //304pi/512
   sin[817]  =  14'b11000000001011;     //305pi/512
   cos[817]  =  14'b00000100101101;     //305pi/512
   sin[818]  =  14'b11000000001010;     //306pi/512
   cos[818]  =  14'b00000100011001;     //306pi/512
   sin[819]  =  14'b11000000001000;     //307pi/512
   cos[819]  =  14'b00000100000101;     //307pi/512
   sin[820]  =  14'b11000000000111;     //308pi/512
   cos[820]  =  14'b00000011110001;     //308pi/512
   sin[821]  =  14'b11000000000110;     //309pi/512
   cos[821]  =  14'b00000011011101;     //309pi/512
   sin[822]  =  14'b11000000000101;     //310pi/512
   cos[822]  =  14'b00000011001000;     //310pi/512
   sin[823]  =  14'b11000000000100;     //311pi/512
   cos[823]  =  14'b00000010110100;     //311pi/512
   sin[824]  =  14'b11000000000011;     //312pi/512
   cos[824]  =  14'b00000010100000;     //312pi/512
   sin[825]  =  14'b11000000000010;     //313pi/512
   cos[825]  =  14'b00000010001100;     //313pi/512
   sin[826]  =  14'b11000000000010;     //314pi/512
   cos[826]  =  14'b00000001111000;     //314pi/512
   sin[827]  =  14'b11000000000001;     //315pi/512
   cos[827]  =  14'b00000001100100;     //315pi/512
   sin[828]  =  14'b11000000000001;     //316pi/512
   cos[828]  =  14'b00000001010000;     //316pi/512
   sin[829]  =  14'b11000000000000;     //317pi/512
   cos[829]  =  14'b00000000111100;     //317pi/512
   sin[830]  =  14'b11000000000000;     //318pi/512
   cos[830]  =  14'b00000000101000;     //318pi/512
   sin[831]  =  14'b11000000000000;     //319pi/512
   cos[831]  =  14'b00000000010100;     //319pi/512
   sin[832]  =  14'b11000000000000;     //320pi/512
   cos[832]  =  14'b00000000000000;     //320pi/512
   sin[833]  =  14'b11000000000000;     //321pi/512
   cos[833]  =  14'b11111111101100;     //321pi/512
   sin[834]  =  14'b11000000000000;     //322pi/512
   cos[834]  =  14'b11111111011000;     //322pi/512
   sin[835]  =  14'b11000000000000;     //323pi/512
   cos[835]  =  14'b11111111000100;     //323pi/512
   sin[836]  =  14'b11000000000001;     //324pi/512
   cos[836]  =  14'b11111110110000;     //324pi/512
   sin[837]  =  14'b11000000000001;     //325pi/512
   cos[837]  =  14'b11111110011011;     //325pi/512
   sin[838]  =  14'b11000000000010;     //326pi/512
   cos[838]  =  14'b11111110000111;     //326pi/512
   sin[839]  =  14'b11000000000010;     //327pi/512
   cos[839]  =  14'b11111101110011;     //327pi/512
   sin[840]  =  14'b11000000000011;     //328pi/512
   cos[840]  =  14'b11111101011111;     //328pi/512
   sin[841]  =  14'b11000000000100;     //329pi/512
   cos[841]  =  14'b11111101001011;     //329pi/512
   sin[842]  =  14'b11000000000101;     //330pi/512
   cos[842]  =  14'b11111100110111;     //330pi/512
   sin[843]  =  14'b11000000000110;     //331pi/512
   cos[843]  =  14'b11111100100011;     //331pi/512
   sin[844]  =  14'b11000000000111;     //332pi/512
   cos[844]  =  14'b11111100001111;     //332pi/512
   sin[845]  =  14'b11000000001000;     //333pi/512
   cos[845]  =  14'b11111011111011;     //333pi/512
   sin[846]  =  14'b11000000001010;     //334pi/512
   cos[846]  =  14'b11111011100111;     //334pi/512
   sin[847]  =  14'b11000000001011;     //335pi/512
   cos[847]  =  14'b11111011010011;     //335pi/512
   sin[848]  =  14'b11000000001101;     //336pi/512
   cos[848]  =  14'b11111010111111;     //336pi/512
   sin[849]  =  14'b11000000001110;     //337pi/512
   cos[849]  =  14'b11111010101011;     //337pi/512
   sin[850]  =  14'b11000000010000;     //338pi/512
   cos[850]  =  14'b11111010010111;     //338pi/512
   sin[851]  =  14'b11000000010010;     //339pi/512
   cos[851]  =  14'b11111010000011;     //339pi/512
   sin[852]  =  14'b11000000010100;     //340pi/512
   cos[852]  =  14'b11111001101111;     //340pi/512
   sin[853]  =  14'b11000000010110;     //341pi/512
   cos[853]  =  14'b11111001011011;     //341pi/512
   sin[854]  =  14'b11000000011000;     //342pi/512
   cos[854]  =  14'b11111001000111;     //342pi/512
   sin[855]  =  14'b11000000011010;     //343pi/512
   cos[855]  =  14'b11111000110011;     //343pi/512
   sin[856]  =  14'b11000000011100;     //344pi/512
   cos[856]  =  14'b11111000011111;     //344pi/512
   sin[857]  =  14'b11000000011111;     //345pi/512
   cos[857]  =  14'b11111000001011;     //345pi/512
   sin[858]  =  14'b11000000100001;     //346pi/512
   cos[858]  =  14'b11110111110111;     //346pi/512
   sin[859]  =  14'b11000000100100;     //347pi/512
   cos[859]  =  14'b11110111100011;     //347pi/512
   sin[860]  =  14'b11000000100111;     //348pi/512
   cos[860]  =  14'b11110111001111;     //348pi/512
   sin[861]  =  14'b11000000101001;     //349pi/512
   cos[861]  =  14'b11110110111011;     //349pi/512
   sin[862]  =  14'b11000000101100;     //350pi/512
   cos[862]  =  14'b11110110100111;     //350pi/512
   sin[863]  =  14'b11000000101111;     //351pi/512
   cos[863]  =  14'b11110110010011;     //351pi/512
   sin[864]  =  14'b11000000110010;     //352pi/512
   cos[864]  =  14'b11110101111111;     //352pi/512
   sin[865]  =  14'b11000000110110;     //353pi/512
   cos[865]  =  14'b11110101101011;     //353pi/512
   sin[866]  =  14'b11000000111001;     //354pi/512
   cos[866]  =  14'b11110101011000;     //354pi/512
   sin[867]  =  14'b11000000111100;     //355pi/512
   cos[867]  =  14'b11110101000100;     //355pi/512
   sin[868]  =  14'b11000001000000;     //356pi/512
   cos[868]  =  14'b11110100110000;     //356pi/512
   sin[869]  =  14'b11000001000011;     //357pi/512
   cos[869]  =  14'b11110100011100;     //357pi/512
   sin[870]  =  14'b11000001000111;     //358pi/512
   cos[870]  =  14'b11110100001000;     //358pi/512
   sin[871]  =  14'b11000001001011;     //359pi/512
   cos[871]  =  14'b11110011110101;     //359pi/512
   sin[872]  =  14'b11000001001111;     //360pi/512
   cos[872]  =  14'b11110011100001;     //360pi/512
   sin[873]  =  14'b11000001010011;     //361pi/512
   cos[873]  =  14'b11110011001101;     //361pi/512
   sin[874]  =  14'b11000001010111;     //362pi/512
   cos[874]  =  14'b11110010111010;     //362pi/512
   sin[875]  =  14'b11000001011011;     //363pi/512
   cos[875]  =  14'b11110010100110;     //363pi/512
   sin[876]  =  14'b11000001011111;     //364pi/512
   cos[876]  =  14'b11110010010010;     //364pi/512
   sin[877]  =  14'b11000001100100;     //365pi/512
   cos[877]  =  14'b11110001111111;     //365pi/512
   sin[878]  =  14'b11000001101000;     //366pi/512
   cos[878]  =  14'b11110001101011;     //366pi/512
   sin[879]  =  14'b11000001101101;     //367pi/512
   cos[879]  =  14'b11110001010111;     //367pi/512
   sin[880]  =  14'b11000001110001;     //368pi/512
   cos[880]  =  14'b11110001000100;     //368pi/512
   sin[881]  =  14'b11000001110110;     //369pi/512
   cos[881]  =  14'b11110000110000;     //369pi/512
   sin[882]  =  14'b11000001111011;     //370pi/512
   cos[882]  =  14'b11110000011101;     //370pi/512
   sin[883]  =  14'b11000010000000;     //371pi/512
   cos[883]  =  14'b11110000001001;     //371pi/512
   sin[884]  =  14'b11000010000101;     //372pi/512
   cos[884]  =  14'b11101111110110;     //372pi/512
   sin[885]  =  14'b11000010001010;     //373pi/512
   cos[885]  =  14'b11101111100010;     //373pi/512
   sin[886]  =  14'b11000010001111;     //374pi/512
   cos[886]  =  14'b11101111001111;     //374pi/512
   sin[887]  =  14'b11000010010100;     //375pi/512
   cos[887]  =  14'b11101110111100;     //375pi/512
   sin[888]  =  14'b11000010011010;     //376pi/512
   cos[888]  =  14'b11101110101000;     //376pi/512
   sin[889]  =  14'b11000010011111;     //377pi/512
   cos[889]  =  14'b11101110010101;     //377pi/512
   sin[890]  =  14'b11000010100101;     //378pi/512
   cos[890]  =  14'b11101110000010;     //378pi/512
   sin[891]  =  14'b11000010101011;     //379pi/512
   cos[891]  =  14'b11101101101110;     //379pi/512
   sin[892]  =  14'b11000010110000;     //380pi/512
   cos[892]  =  14'b11101101011011;     //380pi/512
   sin[893]  =  14'b11000010110110;     //381pi/512
   cos[893]  =  14'b11101101001000;     //381pi/512
   sin[894]  =  14'b11000010111100;     //382pi/512
   cos[894]  =  14'b11101100110101;     //382pi/512
   sin[895]  =  14'b11000011000010;     //383pi/512
   cos[895]  =  14'b11101100100001;     //383pi/512
   sin[896]  =  14'b11000011001000;     //384pi/512
   cos[896]  =  14'b11101100001110;     //384pi/512
   sin[897]  =  14'b11000011001111;     //385pi/512
   cos[897]  =  14'b11101011111011;     //385pi/512
   sin[898]  =  14'b11000011010101;     //386pi/512
   cos[898]  =  14'b11101011101000;     //386pi/512
   sin[899]  =  14'b11000011011100;     //387pi/512
   cos[899]  =  14'b11101011010101;     //387pi/512
   sin[900]  =  14'b11000011100010;     //388pi/512
   cos[900]  =  14'b11101011000010;     //388pi/512
   sin[901]  =  14'b11000011101001;     //389pi/512
   cos[901]  =  14'b11101010101111;     //389pi/512
   sin[902]  =  14'b11000011101111;     //390pi/512
   cos[902]  =  14'b11101010011100;     //390pi/512
   sin[903]  =  14'b11000011110110;     //391pi/512
   cos[903]  =  14'b11101010001001;     //391pi/512
   sin[904]  =  14'b11000011111101;     //392pi/512
   cos[904]  =  14'b11101001110110;     //392pi/512
   sin[905]  =  14'b11000100000100;     //393pi/512
   cos[905]  =  14'b11101001100011;     //393pi/512
   sin[906]  =  14'b11000100001011;     //394pi/512
   cos[906]  =  14'b11101001010001;     //394pi/512
   sin[907]  =  14'b11000100010010;     //395pi/512
   cos[907]  =  14'b11101000111110;     //395pi/512
   sin[908]  =  14'b11000100011010;     //396pi/512
   cos[908]  =  14'b11101000101011;     //396pi/512
   sin[909]  =  14'b11000100100001;     //397pi/512
   cos[909]  =  14'b11101000011000;     //397pi/512
   sin[910]  =  14'b11000100101001;     //398pi/512
   cos[910]  =  14'b11101000000110;     //398pi/512
   sin[911]  =  14'b11000100110000;     //399pi/512
   cos[911]  =  14'b11100111110011;     //399pi/512
   sin[912]  =  14'b11000100111000;     //400pi/512
   cos[912]  =  14'b11100111100001;     //400pi/512
   sin[913]  =  14'b11000101000000;     //401pi/512
   cos[913]  =  14'b11100111001110;     //401pi/512
   sin[914]  =  14'b11000101000111;     //402pi/512
   cos[914]  =  14'b11100110111011;     //402pi/512
   sin[915]  =  14'b11000101001111;     //403pi/512
   cos[915]  =  14'b11100110101001;     //403pi/512
   sin[916]  =  14'b11000101010111;     //404pi/512
   cos[916]  =  14'b11100110010111;     //404pi/512
   sin[917]  =  14'b11000101011111;     //405pi/512
   cos[917]  =  14'b11100110000100;     //405pi/512
   sin[918]  =  14'b11000101101000;     //406pi/512
   cos[918]  =  14'b11100101110010;     //406pi/512
   sin[919]  =  14'b11000101110000;     //407pi/512
   cos[919]  =  14'b11100101011111;     //407pi/512
   sin[920]  =  14'b11000101111000;     //408pi/512
   cos[920]  =  14'b11100101001101;     //408pi/512
   sin[921]  =  14'b11000110000001;     //409pi/512
   cos[921]  =  14'b11100100111011;     //409pi/512
   sin[922]  =  14'b11000110001001;     //410pi/512
   cos[922]  =  14'b11100100101001;     //410pi/512
   sin[923]  =  14'b11000110010010;     //411pi/512
   cos[923]  =  14'b11100100010111;     //411pi/512
   sin[924]  =  14'b11000110011011;     //412pi/512
   cos[924]  =  14'b11100100000100;     //412pi/512
   sin[925]  =  14'b11000110100011;     //413pi/512
   cos[925]  =  14'b11100011110010;     //413pi/512
   sin[926]  =  14'b11000110101100;     //414pi/512
   cos[926]  =  14'b11100011100000;     //414pi/512
   sin[927]  =  14'b11000110110101;     //415pi/512
   cos[927]  =  14'b11100011001110;     //415pi/512
   sin[928]  =  14'b11000110111110;     //416pi/512
   cos[928]  =  14'b11100010111100;     //416pi/512
   sin[929]  =  14'b11000111001000;     //417pi/512
   cos[929]  =  14'b11100010101011;     //417pi/512
   sin[930]  =  14'b11000111010001;     //418pi/512
   cos[930]  =  14'b11100010011001;     //418pi/512
   sin[931]  =  14'b11000111011010;     //419pi/512
   cos[931]  =  14'b11100010000111;     //419pi/512
   sin[932]  =  14'b11000111100100;     //420pi/512
   cos[932]  =  14'b11100001110101;     //420pi/512
   sin[933]  =  14'b11000111101101;     //421pi/512
   cos[933]  =  14'b11100001100011;     //421pi/512
   sin[934]  =  14'b11000111110111;     //422pi/512
   cos[934]  =  14'b11100001010010;     //422pi/512
   sin[935]  =  14'b11001000000000;     //423pi/512
   cos[935]  =  14'b11100001000000;     //423pi/512
   sin[936]  =  14'b11001000001010;     //424pi/512
   cos[936]  =  14'b11100000101111;     //424pi/512
   sin[937]  =  14'b11001000010100;     //425pi/512
   cos[937]  =  14'b11100000011101;     //425pi/512
   sin[938]  =  14'b11001000011110;     //426pi/512
   cos[938]  =  14'b11100000001100;     //426pi/512
   sin[939]  =  14'b11001000101000;     //427pi/512
   cos[939]  =  14'b11011111111010;     //427pi/512
   sin[940]  =  14'b11001000110010;     //428pi/512
   cos[940]  =  14'b11011111101001;     //428pi/512
   sin[941]  =  14'b11001000111100;     //429pi/512
   cos[941]  =  14'b11011111011000;     //429pi/512
   sin[942]  =  14'b11001001000111;     //430pi/512
   cos[942]  =  14'b11011111000110;     //430pi/512
   sin[943]  =  14'b11001001010001;     //431pi/512
   cos[943]  =  14'b11011110110101;     //431pi/512
   sin[944]  =  14'b11001001011100;     //432pi/512
   cos[944]  =  14'b11011110100100;     //432pi/512
   sin[945]  =  14'b11001001100110;     //433pi/512
   cos[945]  =  14'b11011110010011;     //433pi/512
   sin[946]  =  14'b11001001110001;     //434pi/512
   cos[946]  =  14'b11011110000010;     //434pi/512
   sin[947]  =  14'b11001001111011;     //435pi/512
   cos[947]  =  14'b11011101110001;     //435pi/512
   sin[948]  =  14'b11001010000110;     //436pi/512
   cos[948]  =  14'b11011101100000;     //436pi/512
   sin[949]  =  14'b11001010010001;     //437pi/512
   cos[949]  =  14'b11011101001111;     //437pi/512
   sin[950]  =  14'b11001010011100;     //438pi/512
   cos[950]  =  14'b11011100111110;     //438pi/512
   sin[951]  =  14'b11001010100111;     //439pi/512
   cos[951]  =  14'b11011100101101;     //439pi/512
   sin[952]  =  14'b11001010110010;     //440pi/512
   cos[952]  =  14'b11011100011100;     //440pi/512
   sin[953]  =  14'b11001010111110;     //441pi/512
   cos[953]  =  14'b11011100001100;     //441pi/512
   sin[954]  =  14'b11001011001001;     //442pi/512
   cos[954]  =  14'b11011011111011;     //442pi/512
   sin[955]  =  14'b11001011010100;     //443pi/512
   cos[955]  =  14'b11011011101010;     //443pi/512
   sin[956]  =  14'b11001011100000;     //444pi/512
   cos[956]  =  14'b11011011011010;     //444pi/512
   sin[957]  =  14'b11001011101011;     //445pi/512
   cos[957]  =  14'b11011011001001;     //445pi/512
   sin[958]  =  14'b11001011110111;     //446pi/512
   cos[958]  =  14'b11011010111001;     //446pi/512
   sin[959]  =  14'b11001100000010;     //447pi/512
   cos[959]  =  14'b11011010101001;     //447pi/512
   sin[960]  =  14'b11001100001110;     //448pi/512
   cos[960]  =  14'b11011010011000;     //448pi/512
   sin[961]  =  14'b11001100011010;     //449pi/512
   cos[961]  =  14'b11011010001000;     //449pi/512
   sin[962]  =  14'b11001100100110;     //450pi/512
   cos[962]  =  14'b11011001111000;     //450pi/512
   sin[963]  =  14'b11001100110010;     //451pi/512
   cos[963]  =  14'b11011001101000;     //451pi/512
   sin[964]  =  14'b11001100111110;     //452pi/512
   cos[964]  =  14'b11011001011000;     //452pi/512
   sin[965]  =  14'b11001101001010;     //453pi/512
   cos[965]  =  14'b11011001001000;     //453pi/512
   sin[966]  =  14'b11001101010111;     //454pi/512
   cos[966]  =  14'b11011000111000;     //454pi/512
   sin[967]  =  14'b11001101100011;     //455pi/512
   cos[967]  =  14'b11011000101000;     //455pi/512
   sin[968]  =  14'b11001101101111;     //456pi/512
   cos[968]  =  14'b11011000011000;     //456pi/512
   sin[969]  =  14'b11001101111100;     //457pi/512
   cos[969]  =  14'b11011000001000;     //457pi/512
   sin[970]  =  14'b11001110001000;     //458pi/512
   cos[970]  =  14'b11010111111001;     //458pi/512
   sin[971]  =  14'b11001110010101;     //459pi/512
   cos[971]  =  14'b11010111101001;     //459pi/512
   sin[972]  =  14'b11001110100010;     //460pi/512
   cos[972]  =  14'b11010111011010;     //460pi/512
   sin[973]  =  14'b11001110101111;     //461pi/512
   cos[973]  =  14'b11010111001010;     //461pi/512
   sin[974]  =  14'b11001110111011;     //462pi/512
   cos[974]  =  14'b11010110111011;     //462pi/512
   sin[975]  =  14'b11001111001000;     //463pi/512
   cos[975]  =  14'b11010110101011;     //463pi/512
   sin[976]  =  14'b11001111010101;     //464pi/512
   cos[976]  =  14'b11010110011100;     //464pi/512
   sin[977]  =  14'b11001111100010;     //465pi/512
   cos[977]  =  14'b11010110001101;     //465pi/512
   sin[978]  =  14'b11001111110000;     //466pi/512
   cos[978]  =  14'b11010101111101;     //466pi/512
   sin[979]  =  14'b11001111111101;     //467pi/512
   cos[979]  =  14'b11010101101110;     //467pi/512
   sin[980]  =  14'b11010000001010;     //468pi/512
   cos[980]  =  14'b11010101011111;     //468pi/512
   sin[981]  =  14'b11010000011000;     //469pi/512
   cos[981]  =  14'b11010101010000;     //469pi/512
   sin[982]  =  14'b11010000100101;     //470pi/512
   cos[982]  =  14'b11010101000001;     //470pi/512
   sin[983]  =  14'b11010000110011;     //471pi/512
   cos[983]  =  14'b11010100110010;     //471pi/512
   sin[984]  =  14'b11010001000000;     //472pi/512
   cos[984]  =  14'b11010100100100;     //472pi/512
   sin[985]  =  14'b11010001001110;     //473pi/512
   cos[985]  =  14'b11010100010101;     //473pi/512
   sin[986]  =  14'b11010001011100;     //474pi/512
   cos[986]  =  14'b11010100000110;     //474pi/512
   sin[987]  =  14'b11010001101001;     //475pi/512
   cos[987]  =  14'b11010011111000;     //475pi/512
   sin[988]  =  14'b11010001110111;     //476pi/512
   cos[988]  =  14'b11010011101001;     //476pi/512
   sin[989]  =  14'b11010010000101;     //477pi/512
   cos[989]  =  14'b11010011011011;     //477pi/512
   sin[990]  =  14'b11010010010011;     //478pi/512
   cos[990]  =  14'b11010011001100;     //478pi/512
   sin[991]  =  14'b11010010100010;     //479pi/512
   cos[991]  =  14'b11010010111110;     //479pi/512
   sin[992]  =  14'b11010010110000;     //480pi/512
   cos[992]  =  14'b11010010110000;     //480pi/512
   sin[993]  =  14'b11010010111110;     //481pi/512
   cos[993]  =  14'b11010010100010;     //481pi/512
   sin[994]  =  14'b11010011001100;     //482pi/512
   cos[994]  =  14'b11010010010011;     //482pi/512
   sin[995]  =  14'b11010011011011;     //483pi/512
   cos[995]  =  14'b11010010000101;     //483pi/512
   sin[996]  =  14'b11010011101001;     //484pi/512
   cos[996]  =  14'b11010001110111;     //484pi/512
   sin[997]  =  14'b11010011111000;     //485pi/512
   cos[997]  =  14'b11010001101001;     //485pi/512
   sin[998]  =  14'b11010100000110;     //486pi/512
   cos[998]  =  14'b11010001011100;     //486pi/512
   sin[999]  =  14'b11010100010101;     //487pi/512
   cos[999]  =  14'b11010001001110;     //487pi/512
   sin[1000]  =  14'b11010100100100;     //488pi/512
   cos[1000]  =  14'b11010001000000;     //488pi/512
   sin[1001]  =  14'b11010100110010;     //489pi/512
   cos[1001]  =  14'b11010000110011;     //489pi/512
   sin[1002]  =  14'b11010101000001;     //490pi/512
   cos[1002]  =  14'b11010000100101;     //490pi/512
   sin[1003]  =  14'b11010101010000;     //491pi/512
   cos[1003]  =  14'b11010000011000;     //491pi/512
   sin[1004]  =  14'b11010101011111;     //492pi/512
   cos[1004]  =  14'b11010000001010;     //492pi/512
   sin[1005]  =  14'b11010101101110;     //493pi/512
   cos[1005]  =  14'b11001111111101;     //493pi/512
   sin[1006]  =  14'b11010101111101;     //494pi/512
   cos[1006]  =  14'b11001111110000;     //494pi/512
   sin[1007]  =  14'b11010110001101;     //495pi/512
   cos[1007]  =  14'b11001111100010;     //495pi/512
   sin[1008]  =  14'b11010110011100;     //496pi/512
   cos[1008]  =  14'b11001111010101;     //496pi/512
   sin[1009]  =  14'b11010110101011;     //497pi/512
   cos[1009]  =  14'b11001111001000;     //497pi/512
   sin[1010]  =  14'b11010110111011;     //498pi/512
   cos[1010]  =  14'b11001110111011;     //498pi/512
   sin[1011]  =  14'b11010111001010;     //499pi/512
   cos[1011]  =  14'b11001110101111;     //499pi/512
   sin[1012]  =  14'b11010111011010;     //500pi/512
   cos[1012]  =  14'b11001110100010;     //500pi/512
   sin[1013]  =  14'b11010111101001;     //501pi/512
   cos[1013]  =  14'b11001110010101;     //501pi/512
   sin[1014]  =  14'b11010111111001;     //502pi/512
   cos[1014]  =  14'b11001110001000;     //502pi/512
   sin[1015]  =  14'b11011000001000;     //503pi/512
   cos[1015]  =  14'b11001101111100;     //503pi/512
   sin[1016]  =  14'b11011000011000;     //504pi/512
   cos[1016]  =  14'b11001101101111;     //504pi/512
   sin[1017]  =  14'b11011000101000;     //505pi/512
   cos[1017]  =  14'b11001101100011;     //505pi/512
   sin[1018]  =  14'b11011000111000;     //506pi/512
   cos[1018]  =  14'b11001101010111;     //506pi/512
   sin[1019]  =  14'b11011001001000;     //507pi/512
   cos[1019]  =  14'b11001101001010;     //507pi/512
   sin[1020]  =  14'b11011001011000;     //508pi/512
   cos[1020]  =  14'b11001100111110;     //508pi/512
   sin[1021]  =  14'b11011001101000;     //509pi/512
   cos[1021]  =  14'b11001100110010;     //509pi/512
   sin[1022]  =  14'b11011001111000;     //510pi/512
   cos[1022]  =  14'b11001100100110;     //510pi/512
   sin[1023]  =  14'b11011010001000;     //511pi/512
   cos[1023]  =  14'b11001100011010;     //511pi/512
end
endmodule