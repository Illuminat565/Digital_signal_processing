
module  TWIDLE_16_bit  (
    input   [10:0]   rd_ptr_angle,

    output  signed [15:0]   cos_data,
    output  signed [15:0]   sin_data
 );

wire signed [15:0]  cos  [511:0];
wire signed [15:0]  sin  [511:0];

assign cos_data =    cos [rd_ptr_angle];
assign sin_data =    sin [rd_ptr_angle];

  assign sin[0]  =  16'b0000_0000_0000_0000;     //0pi/512
  assign cos[0]  =  16'b0100_0000_0000_0000;     //0pi/512
  assign sin[1]  =  16'b1111_1111_1001_1011;     //1pi/512
  assign cos[1]  =  16'b0011_1111_1111_1111;     //1pi/512
  assign sin[2]  =  16'b1111_1111_0011_0111;     //2pi/512
  assign cos[2]  =  16'b0011_1111_1111_1110;     //2pi/512
  assign sin[3]  =  16'b1111_1110_1101_0010;     //3pi/512
  assign cos[3]  =  16'b0011_1111_1111_1101;     //3pi/512
  assign sin[4]  =  16'b1111_1110_0110_1110;     //4pi/512
  assign cos[4]  =  16'b0011_1111_1111_1011;     //4pi/512
  assign sin[5]  =  16'b1111_1110_0000_1001;     //5pi/512
  assign cos[5]  =  16'b0011_1111_1111_1000;     //5pi/512
  assign sin[6]  =  16'b1111_1101_1010_0101;     //6pi/512
  assign cos[6]  =  16'b0011_1111_1111_0100;     //6pi/512
  assign sin[7]  =  16'b1111_1101_0100_0000;     //7pi/512
  assign cos[7]  =  16'b0011_1111_1111_0000;     //7pi/512
  assign sin[8]  =  16'b1111_1100_1101_1100;     //8pi/512
  assign cos[8]  =  16'b0011_1111_1110_1100;     //8pi/512
  assign sin[9]  =  16'b1111_1100_0111_1000;     //9pi/512
  assign cos[9]  =  16'b0011_1111_1110_0111;     //9pi/512
  assign sin[10]  =  16'b1111_1100_0001_0011;     //10pi/512
  assign cos[10]  =  16'b0011_1111_1110_0001;     //10pi/512
  assign sin[11]  =  16'b1111_1011_1010_1111;     //11pi/512
  assign cos[11]  =  16'b0011_1111_1101_1010;     //11pi/512
  assign sin[12]  =  16'b1111_1011_0100_1011;     //12pi/512
  assign cos[12]  =  16'b0011_1111_1101_0011;     //12pi/512
  assign sin[13]  =  16'b1111_1010_1110_0110;     //13pi/512
  assign cos[13]  =  16'b0011_1111_1100_1011;     //13pi/512
  assign sin[14]  =  16'b1111_1010_1000_0010;     //14pi/512
  assign cos[14]  =  16'b0011_1111_1100_0011;     //14pi/512
  assign sin[15]  =  16'b1111_1010_0001_1110;     //15pi/512
  assign cos[15]  =  16'b0011_1111_1011_1010;     //15pi/512
  assign sin[16]  =  16'b1111_1001_1011_1010;     //16pi/512
  assign cos[16]  =  16'b0011_1111_1011_0001;     //16pi/512
  assign sin[17]  =  16'b1111_1001_0101_0110;     //17pi/512
  assign cos[17]  =  16'b0011_1111_1010_0110;     //17pi/512
  assign sin[18]  =  16'b1111_1000_1111_0010;     //18pi/512
  assign cos[18]  =  16'b0011_1111_1001_1100;     //18pi/512
  assign sin[19]  =  16'b1111_1000_1000_1110;     //19pi/512
  assign cos[19]  =  16'b0011_1111_1001_0000;     //19pi/512
  assign sin[20]  =  16'b1111_1000_0010_1010;     //20pi/512
  assign cos[20]  =  16'b0011_1111_1000_0100;     //20pi/512
  assign sin[21]  =  16'b1111_0111_1100_0111;     //21pi/512
  assign cos[21]  =  16'b0011_1111_0111_1000;     //21pi/512
  assign sin[22]  =  16'b1111_0111_0110_0011;     //22pi/512
  assign cos[22]  =  16'b0011_1111_0110_1010;     //22pi/512
  assign sin[23]  =  16'b1111_0110_1111_1111;     //23pi/512
  assign cos[23]  =  16'b0011_1111_0101_1101;     //23pi/512
  assign sin[24]  =  16'b1111_0110_1001_1100;     //24pi/512
  assign cos[24]  =  16'b0011_1111_0100_1110;     //24pi/512
  assign sin[25]  =  16'b1111_0110_0011_1001;     //25pi/512
  assign cos[25]  =  16'b0011_1111_0011_1111;     //25pi/512
  assign sin[26]  =  16'b1111_0101_1101_0101;     //26pi/512
  assign cos[26]  =  16'b0011_1111_0010_1111;     //26pi/512
  assign sin[27]  =  16'b1111_0101_0111_0010;     //27pi/512
  assign cos[27]  =  16'b0011_1111_0001_1111;     //27pi/512
  assign sin[28]  =  16'b1111_0101_0000_1111;     //28pi/512
  assign cos[28]  =  16'b0011_1111_0000_1110;     //28pi/512
  assign sin[29]  =  16'b1111_0100_1010_1100;     //29pi/512
  assign cos[29]  =  16'b0011_1110_1111_1101;     //29pi/512
  assign sin[30]  =  16'b1111_0100_0100_1001;     //30pi/512
  assign cos[30]  =  16'b0011_1110_1110_1011;     //30pi/512
  assign sin[31]  =  16'b1111_0011_1110_0110;     //31pi/512
  assign cos[31]  =  16'b0011_1110_1101_1000;     //31pi/512
  assign sin[32]  =  16'b1111_0011_1000_0100;     //32pi/512
  assign cos[32]  =  16'b0011_1110_1100_0101;     //32pi/512
  assign sin[33]  =  16'b1111_0011_0010_0001;     //33pi/512
  assign cos[33]  =  16'b0011_1110_1011_0001;     //33pi/512
  assign sin[34]  =  16'b1111_0010_1011_1111;     //34pi/512
  assign cos[34]  =  16'b0011_1110_1001_1100;     //34pi/512
  assign sin[35]  =  16'b1111_0010_0101_1100;     //35pi/512
  assign cos[35]  =  16'b0011_1110_1000_0111;     //35pi/512
  assign sin[36]  =  16'b1111_0001_1111_1010;     //36pi/512
  assign cos[36]  =  16'b0011_1110_0111_0001;     //36pi/512
  assign sin[37]  =  16'b1111_0001_1001_1000;     //37pi/512
  assign cos[37]  =  16'b0011_1110_0101_1011;     //37pi/512
  assign sin[38]  =  16'b1111_0001_0011_0110;     //38pi/512
  assign cos[38]  =  16'b0011_1110_0100_0100;     //38pi/512
  assign sin[39]  =  16'b1111_0000_1101_0101;     //39pi/512
  assign cos[39]  =  16'b0011_1110_0010_1101;     //39pi/512
  assign sin[40]  =  16'b1111_0000_0111_0011;     //40pi/512
  assign cos[40]  =  16'b0011_1110_0001_0100;     //40pi/512
  assign sin[41]  =  16'b1111_0000_0001_0010;     //41pi/512
  assign cos[41]  =  16'b0011_1101_1111_1100;     //41pi/512
  assign sin[42]  =  16'b1110_1111_1011_0000;     //42pi/512
  assign cos[42]  =  16'b0011_1101_1110_0010;     //42pi/512
  assign sin[43]  =  16'b1110_1111_0100_1111;     //43pi/512
  assign cos[43]  =  16'b0011_1101_1100_1001;     //43pi/512
  assign sin[44]  =  16'b1110_1110_1110_1110;     //44pi/512
  assign cos[44]  =  16'b0011_1101_1010_1110;     //44pi/512
  assign sin[45]  =  16'b1110_1110_1000_1101;     //45pi/512
  assign cos[45]  =  16'b0011_1101_1001_0011;     //45pi/512
  assign sin[46]  =  16'b1110_1110_0010_1101;     //46pi/512
  assign cos[46]  =  16'b0011_1101_0111_0111;     //46pi/512
  assign sin[47]  =  16'b1110_1101_1100_1100;     //47pi/512
  assign cos[47]  =  16'b0011_1101_0101_1011;     //47pi/512
  assign sin[48]  =  16'b1110_1101_0110_1100;     //48pi/512
  assign cos[48]  =  16'b0011_1101_0011_1110;     //48pi/512
  assign sin[49]  =  16'b1110_1101_0000_1100;     //49pi/512
  assign cos[49]  =  16'b0011_1101_0010_0001;     //49pi/512
  assign sin[50]  =  16'b1110_1100_1010_1100;     //50pi/512
  assign cos[50]  =  16'b0011_1101_0000_0010;     //50pi/512
  assign sin[51]  =  16'b1110_1100_0100_1100;     //51pi/512
  assign cos[51]  =  16'b0011_1100_1110_0100;     //51pi/512
  assign sin[52]  =  16'b1110_1011_1110_1101;     //52pi/512
  assign cos[52]  =  16'b0011_1100_1100_0101;     //52pi/512
  assign sin[53]  =  16'b1110_1011_1000_1101;     //53pi/512
  assign cos[53]  =  16'b0011_1100_1010_0101;     //53pi/512
  assign sin[54]  =  16'b1110_1011_0010_1110;     //54pi/512
  assign cos[54]  =  16'b0011_1100_1000_0100;     //54pi/512
  assign sin[55]  =  16'b1110_1010_1100_1111;     //55pi/512
  assign cos[55]  =  16'b0011_1100_0110_0011;     //55pi/512
  assign sin[56]  =  16'b1110_1010_0111_0000;     //56pi/512
  assign cos[56]  =  16'b0011_1100_0100_0010;     //56pi/512
  assign sin[57]  =  16'b1110_1010_0001_0010;     //57pi/512
  assign cos[57]  =  16'b0011_1100_0010_0000;     //57pi/512
  assign sin[58]  =  16'b1110_1001_1011_0100;     //58pi/512
  assign cos[58]  =  16'b0011_1011_1111_1101;     //58pi/512
  assign sin[59]  =  16'b1110_1001_0101_0101;     //59pi/512
  assign cos[59]  =  16'b0011_1011_1101_1010;     //59pi/512
  assign sin[60]  =  16'b1110_1000_1111_0111;     //60pi/512
  assign cos[60]  =  16'b0011_1011_1011_0110;     //60pi/512
  assign sin[61]  =  16'b1110_1000_1001_1010;     //61pi/512
  assign cos[61]  =  16'b0011_1011_1001_0001;     //61pi/512
  assign sin[62]  =  16'b1110_1000_0011_1100;     //62pi/512
  assign cos[62]  =  16'b0011_1011_0110_1100;     //62pi/512
  assign sin[63]  =  16'b1110_0111_1101_1111;     //63pi/512
  assign cos[63]  =  16'b0011_1011_0100_0111;     //63pi/512
  assign sin[64]  =  16'b1110_0111_1000_0010;     //64pi/512
  assign cos[64]  =  16'b0011_1011_0010_0000;     //64pi/512
  assign sin[65]  =  16'b1110_0111_0010_0101;     //65pi/512
  assign cos[65]  =  16'b0011_1010_1111_1010;     //65pi/512
  assign sin[66]  =  16'b1110_0110_1100_1001;     //66pi/512
  assign cos[66]  =  16'b0011_1010_1101_0010;     //66pi/512
  assign sin[67]  =  16'b1110_0110_0110_1101;     //67pi/512
  assign cos[67]  =  16'b0011_1010_1010_1010;     //67pi/512
  assign sin[68]  =  16'b1110_0110_0001_0001;     //68pi/512
  assign cos[68]  =  16'b0011_1010_1000_0010;     //68pi/512
  assign sin[69]  =  16'b1110_0101_1011_0101;     //69pi/512
  assign cos[69]  =  16'b0011_1010_0101_1001;     //69pi/512
  assign sin[70]  =  16'b1110_0101_0101_1001;     //70pi/512
  assign cos[70]  =  16'b0011_1010_0010_1111;     //70pi/512
  assign sin[71]  =  16'b1110_0100_1111_1110;     //71pi/512
  assign cos[71]  =  16'b0011_1010_0000_0101;     //71pi/512
  assign sin[72]  =  16'b1110_0100_1010_0011;     //72pi/512
  assign cos[72]  =  16'b0011_1001_1101_1010;     //72pi/512
  assign sin[73]  =  16'b1110_0100_0100_1000;     //73pi/512
  assign cos[73]  =  16'b0011_1001_1010_1111;     //73pi/512
  assign sin[74]  =  16'b1110_0011_1110_1110;     //74pi/512
  assign cos[74]  =  16'b0011_1001_1000_0011;     //74pi/512
  assign sin[75]  =  16'b1110_0011_1001_0100;     //75pi/512
  assign cos[75]  =  16'b0011_1001_0101_0111;     //75pi/512
  assign sin[76]  =  16'b1110_0011_0011_1010;     //76pi/512
  assign cos[76]  =  16'b0011_1001_0010_1010;     //76pi/512
  assign sin[77]  =  16'b1110_0010_1110_0000;     //77pi/512
  assign cos[77]  =  16'b0011_1000_1111_1101;     //77pi/512
  assign sin[78]  =  16'b1110_0010_1000_0111;     //78pi/512
  assign cos[78]  =  16'b0011_1000_1100_1111;     //78pi/512
  assign sin[79]  =  16'b1110_0010_0010_1101;     //79pi/512
  assign cos[79]  =  16'b0011_1000_1010_0000;     //79pi/512
  assign sin[80]  =  16'b1110_0001_1101_0101;     //80pi/512
  assign cos[80]  =  16'b0011_1000_0111_0001;     //80pi/512
  assign sin[81]  =  16'b1110_0001_0111_1100;     //81pi/512
  assign cos[81]  =  16'b0011_1000_0100_0001;     //81pi/512
  assign sin[82]  =  16'b1110_0001_0010_0100;     //82pi/512
  assign cos[82]  =  16'b0011_1000_0001_0001;     //82pi/512
  assign sin[83]  =  16'b1110_0000_1100_1100;     //83pi/512
  assign cos[83]  =  16'b0011_0111_1110_0000;     //83pi/512
  assign sin[84]  =  16'b1110_0000_0111_0100;     //84pi/512
  assign cos[84]  =  16'b0011_0111_1010_1111;     //84pi/512
  assign sin[85]  =  16'b1110_0000_0001_1101;     //85pi/512
  assign cos[85]  =  16'b0011_0111_0111_1101;     //85pi/512
  assign sin[86]  =  16'b1101_1111_1100_0110;     //86pi/512
  assign cos[86]  =  16'b0011_0111_0100_1011;     //86pi/512
  assign sin[87]  =  16'b1101_1111_0110_1111;     //87pi/512
  assign cos[87]  =  16'b0011_0111_0001_1000;     //87pi/512
  assign sin[88]  =  16'b1101_1111_0001_1001;     //88pi/512
  assign cos[88]  =  16'b0011_0110_1110_0101;     //88pi/512
  assign sin[89]  =  16'b1101_1110_1100_0011;     //89pi/512
  assign cos[89]  =  16'b0011_0110_1011_0001;     //89pi/512
  assign sin[90]  =  16'b1101_1110_0110_1101;     //90pi/512
  assign cos[90]  =  16'b0011_0110_0111_1100;     //90pi/512
  assign sin[91]  =  16'b1101_1110_0001_1000;     //91pi/512
  assign cos[91]  =  16'b0011_0110_0100_0111;     //91pi/512
  assign sin[92]  =  16'b1101_1101_1100_0011;     //92pi/512
  assign cos[92]  =  16'b0011_0110_0001_0010;     //92pi/512
  assign sin[93]  =  16'b1101_1101_0110_1110;     //93pi/512
  assign cos[93]  =  16'b0011_0101_1101_1100;     //93pi/512
  assign sin[94]  =  16'b1101_1101_0001_1001;     //94pi/512
  assign cos[94]  =  16'b0011_0101_1010_0101;     //94pi/512
  assign sin[95]  =  16'b1101_1100_1100_0101;     //95pi/512
  assign cos[95]  =  16'b0011_0101_0110_1110;     //95pi/512
  assign sin[96]  =  16'b1101_1100_0111_0010;     //96pi/512
  assign cos[96]  =  16'b0011_0101_0011_0110;     //96pi/512
  assign sin[97]  =  16'b1101_1100_0001_1110;     //97pi/512
  assign cos[97]  =  16'b0011_0100_1111_1110;     //97pi/512
  assign sin[98]  =  16'b1101_1011_1100_1011;     //98pi/512
  assign cos[98]  =  16'b0011_0100_1100_0110;     //98pi/512
  assign sin[99]  =  16'b1101_1011_0111_1000;     //99pi/512
  assign cos[99]  =  16'b0011_0100_1000_1100;     //99pi/512
  assign sin[100]  =  16'b1101_1011_0010_0110;     //100pi/512
  assign cos[100]  =  16'b0011_0100_0101_0011;     //100pi/512
  assign sin[101]  =  16'b1101_1010_1101_0100;     //101pi/512
  assign cos[101]  =  16'b0011_0100_0001_1001;     //101pi/512
  assign sin[102]  =  16'b1101_1010_1000_0010;     //102pi/512
  assign cos[102]  =  16'b0011_0011_1101_1110;     //102pi/512
  assign sin[103]  =  16'b1101_1010_0011_0001;     //103pi/512
  assign cos[103]  =  16'b0011_0011_1010_0011;     //103pi/512
  assign sin[104]  =  16'b1101_1001_1110_0000;     //104pi/512
  assign cos[104]  =  16'b0011_0011_0110_0111;     //104pi/512
  assign sin[105]  =  16'b1101_1001_1000_1111;     //105pi/512
  assign cos[105]  =  16'b0011_0011_0010_1011;     //105pi/512
  assign sin[106]  =  16'b1101_1001_0011_1111;     //106pi/512
  assign cos[106]  =  16'b0011_0010_1110_1110;     //106pi/512
  assign sin[107]  =  16'b1101_1000_1110_1111;     //107pi/512
  assign cos[107]  =  16'b0011_0010_1011_0001;     //107pi/512
  assign sin[108]  =  16'b1101_1000_1010_0000;     //108pi/512
  assign cos[108]  =  16'b0011_0010_0111_0100;     //108pi/512
  assign sin[109]  =  16'b1101_1000_0101_0001;     //109pi/512
  assign cos[109]  =  16'b0011_0010_0011_0110;     //109pi/512
  assign sin[110]  =  16'b1101_1000_0000_0010;     //110pi/512
  assign cos[110]  =  16'b0011_0001_1111_0111;     //110pi/512
  assign sin[111]  =  16'b1101_0111_1011_0100;     //111pi/512
  assign cos[111]  =  16'b0011_0001_1011_1000;     //111pi/512
  assign sin[112]  =  16'b1101_0111_0110_0110;     //112pi/512
  assign cos[112]  =  16'b0011_0001_0111_1001;     //112pi/512
  assign sin[113]  =  16'b1101_0111_0001_1001;     //113pi/512
  assign cos[113]  =  16'b0011_0001_0011_1000;     //113pi/512
  assign sin[114]  =  16'b1101_0110_1100_1011;     //114pi/512
  assign cos[114]  =  16'b0011_0000_1111_1000;     //114pi/512
  assign sin[115]  =  16'b1101_0110_0111_1111;     //115pi/512
  assign cos[115]  =  16'b0011_0000_1011_0111;     //115pi/512
  assign sin[116]  =  16'b1101_0110_0011_0010;     //116pi/512
  assign cos[116]  =  16'b0011_0000_0111_0110;     //116pi/512
  assign sin[117]  =  16'b1101_0101_1110_0110;     //117pi/512
  assign cos[117]  =  16'b0011_0000_0011_0100;     //117pi/512
  assign sin[118]  =  16'b1101_0101_1001_1011;     //118pi/512
  assign cos[118]  =  16'b0010_1111_1111_0001;     //118pi/512
  assign sin[119]  =  16'b1101_0101_0101_0000;     //119pi/512
  assign cos[119]  =  16'b0010_1111_1010_1111;     //119pi/512
  assign sin[120]  =  16'b1101_0101_0000_0101;     //120pi/512
  assign cos[120]  =  16'b0010_1111_0110_1011;     //120pi/512
  assign sin[121]  =  16'b1101_0100_1011_1011;     //121pi/512
  assign cos[121]  =  16'b0010_1111_0010_1000;     //121pi/512
  assign sin[122]  =  16'b1101_0100_0111_0001;     //122pi/512
  assign cos[122]  =  16'b0010_1110_1110_0011;     //122pi/512
  assign sin[123]  =  16'b1101_0100_0010_1000;     //123pi/512
  assign cos[123]  =  16'b0010_1110_1001_1111;     //123pi/512
  assign sin[124]  =  16'b1101_0011_1101_1111;     //124pi/512
  assign cos[124]  =  16'b0010_1110_0101_1010;     //124pi/512
  assign sin[125]  =  16'b1101_0011_1001_0110;     //125pi/512
  assign cos[125]  =  16'b0010_1110_0001_0100;     //125pi/512
  assign sin[126]  =  16'b1101_0011_0100_1110;     //126pi/512
  assign cos[126]  =  16'b0010_1101_1100_1110;     //126pi/512
  assign sin[127]  =  16'b1101_0011_0000_0110;     //127pi/512
  assign cos[127]  =  16'b0010_1101_1000_1000;     //127pi/512
  assign sin[128]  =  16'b1101_0010_1011_1111;     //128pi/512
  assign cos[128]  =  16'b0010_1101_0100_0001;     //128pi/512
  assign sin[129]  =  16'b1101_0010_0111_1000;     //129pi/512
  assign cos[129]  =  16'b0010_1100_1111_1001;     //129pi/512
  assign sin[130]  =  16'b1101_0010_0011_0001;     //130pi/512
  assign cos[130]  =  16'b0010_1100_1011_0010;     //130pi/512
  assign sin[131]  =  16'b1101_0001_1110_1011;     //131pi/512
  assign cos[131]  =  16'b0010_1100_0110_1010;     //131pi/512
  assign sin[132]  =  16'b1101_0001_1010_0110;     //132pi/512
  assign cos[132]  =  16'b0010_1100_0010_0001;     //132pi/512
  assign sin[133]  =  16'b1101_0001_0110_0001;     //133pi/512
  assign cos[133]  =  16'b0010_1011_1101_1000;     //133pi/512
  assign sin[134]  =  16'b1101_0001_0001_1100;     //134pi/512
  assign cos[134]  =  16'b0010_1011_1000_1110;     //134pi/512
  assign sin[135]  =  16'b1101_0000_1101_1000;     //135pi/512
  assign cos[135]  =  16'b0010_1011_0100_0101;     //135pi/512
  assign sin[136]  =  16'b1101_0000_1001_0100;     //136pi/512
  assign cos[136]  =  16'b0010_1010_1111_1010;     //136pi/512
  assign sin[137]  =  16'b1101_0000_0101_0001;     //137pi/512
  assign cos[137]  =  16'b0010_1010_1011_0000;     //137pi/512
  assign sin[138]  =  16'b1101_0000_0000_1110;     //138pi/512
  assign cos[138]  =  16'b0010_1010_0110_0101;     //138pi/512
  assign sin[139]  =  16'b1100_1111_1100_1100;     //139pi/512
  assign cos[139]  =  16'b0010_1010_0001_1001;     //139pi/512
  assign sin[140]  =  16'b1100_1111_1000_1010;     //140pi/512
  assign cos[140]  =  16'b0010_1001_1100_1101;     //140pi/512
  assign sin[141]  =  16'b1100_1111_0100_1000;     //141pi/512
  assign cos[141]  =  16'b0010_1001_1000_0001;     //141pi/512
  assign sin[142]  =  16'b1100_1111_0000_0111;     //142pi/512
  assign cos[142]  =  16'b0010_1001_0011_0100;     //142pi/512
  assign sin[143]  =  16'b1100_1110_1100_0111;     //143pi/512
  assign cos[143]  =  16'b0010_1000_1110_0111;     //143pi/512
  assign sin[144]  =  16'b1100_1110_1000_0111;     //144pi/512
  assign cos[144]  =  16'b0010_1000_1001_1001;     //144pi/512
  assign sin[145]  =  16'b1100_1110_0100_0111;     //145pi/512
  assign cos[145]  =  16'b0010_1000_0100_1011;     //145pi/512
  assign sin[146]  =  16'b1100_1110_0000_1000;     //146pi/512
  assign cos[146]  =  16'b0010_0111_1111_1101;     //146pi/512
  assign sin[147]  =  16'b1100_1101_1100_1010;     //147pi/512
  assign cos[147]  =  16'b0010_0111_1010_1111;     //147pi/512
  assign sin[148]  =  16'b1100_1101_1000_1100;     //148pi/512
  assign cos[148]  =  16'b0010_0111_0101_1111;     //148pi/512
  assign sin[149]  =  16'b1100_1101_0100_1110;     //149pi/512
  assign cos[149]  =  16'b0010_0111_0001_0000;     //149pi/512
  assign sin[150]  =  16'b1100_1101_0001_0001;     //150pi/512
  assign cos[150]  =  16'b0010_0110_1100_0000;     //150pi/512
  assign sin[151]  =  16'b1100_1100_1101_0100;     //151pi/512
  assign cos[151]  =  16'b0010_0110_0111_0000;     //151pi/512
  assign sin[152]  =  16'b1100_1100_1001_1000;     //152pi/512
  assign cos[152]  =  16'b0010_0110_0001_1111;     //152pi/512
  assign sin[153]  =  16'b1100_1100_0101_1101;     //153pi/512
  assign cos[153]  =  16'b0010_0101_1100_1111;     //153pi/512
  assign sin[154]  =  16'b1100_1100_0010_0001;     //154pi/512
  assign cos[154]  =  16'b0010_0101_0111_1101;     //154pi/512
  assign sin[155]  =  16'b1100_1011_1110_0111;     //155pi/512
  assign cos[155]  =  16'b0010_0101_0010_1100;     //155pi/512
  assign sin[156]  =  16'b1100_1011_1010_1101;     //156pi/512
  assign cos[156]  =  16'b0010_0100_1101_1010;     //156pi/512
  assign sin[157]  =  16'b1100_1011_0111_0011;     //157pi/512
  assign cos[157]  =  16'b0010_0100_1000_0111;     //157pi/512
  assign sin[158]  =  16'b1100_1011_0011_1010;     //158pi/512
  assign cos[158]  =  16'b0010_0100_0011_0100;     //158pi/512
  assign sin[159]  =  16'b1100_1011_0000_0001;     //159pi/512
  assign cos[159]  =  16'b0010_0011_1110_0001;     //159pi/512
  assign sin[160]  =  16'b1100_1010_1100_1001;     //160pi/512
  assign cos[160]  =  16'b0010_0011_1000_1110;     //160pi/512
  assign sin[161]  =  16'b1100_1010_1001_0010;     //161pi/512
  assign cos[161]  =  16'b0010_0011_0011_1010;     //161pi/512
  assign sin[162]  =  16'b1100_1010_0101_1011;     //162pi/512
  assign cos[162]  =  16'b0010_0010_1110_0110;     //162pi/512
  assign sin[163]  =  16'b1100_1010_0010_0100;     //163pi/512
  assign cos[163]  =  16'b0010_0010_1001_0010;     //163pi/512
  assign sin[164]  =  16'b1100_1001_1110_1110;     //164pi/512
  assign cos[164]  =  16'b0010_0010_0011_1101;     //164pi/512
  assign sin[165]  =  16'b1100_1001_1011_1000;     //165pi/512
  assign cos[165]  =  16'b0010_0001_1110_1000;     //165pi/512
  assign sin[166]  =  16'b1100_1001_1000_0011;     //166pi/512
  assign cos[166]  =  16'b0010_0001_1001_0010;     //166pi/512
  assign sin[167]  =  16'b1100_1001_0100_1111;     //167pi/512
  assign cos[167]  =  16'b0010_0001_0011_1101;     //167pi/512
  assign sin[168]  =  16'b1100_1001_0001_1011;     //168pi/512
  assign cos[168]  =  16'b0010_0000_1110_0111;     //168pi/512
  assign sin[169]  =  16'b1100_1000_1110_1000;     //169pi/512
  assign cos[169]  =  16'b0010_0000_1001_0000;     //169pi/512
  assign sin[170]  =  16'b1100_1000_1011_0101;     //170pi/512
  assign cos[170]  =  16'b0010_0000_0011_1001;     //170pi/512
  assign sin[171]  =  16'b1100_1000_1000_0010;     //171pi/512
  assign cos[171]  =  16'b0001_1111_1110_0010;     //171pi/512
  assign sin[172]  =  16'b1100_1000_0101_0000;     //172pi/512
  assign cos[172]  =  16'b0001_1111_1000_1011;     //172pi/512
  assign sin[173]  =  16'b1100_1000_0001_1111;     //173pi/512
  assign cos[173]  =  16'b0001_1111_0011_0100;     //173pi/512
  assign sin[174]  =  16'b1100_0111_1110_1110;     //174pi/512
  assign cos[174]  =  16'b0001_1110_1101_1100;     //174pi/512
  assign sin[175]  =  16'b1100_0111_1011_1110;     //175pi/512
  assign cos[175]  =  16'b0001_1110_1000_0011;     //175pi/512
  assign sin[176]  =  16'b1100_0111_1000_1111;     //176pi/512
  assign cos[176]  =  16'b0001_1110_0010_1011;     //176pi/512
  assign sin[177]  =  16'b1100_0111_0101_1111;     //177pi/512
  assign cos[177]  =  16'b0001_1101_1101_0010;     //177pi/512
  assign sin[178]  =  16'b1100_0111_0011_0001;     //178pi/512
  assign cos[178]  =  16'b0001_1101_0111_1001;     //178pi/512
  assign sin[179]  =  16'b1100_0111_0000_0011;     //179pi/512
  assign cos[179]  =  16'b0001_1101_0010_0000;     //179pi/512
  assign sin[180]  =  16'b1100_0110_1101_0101;     //180pi/512
  assign cos[180]  =  16'b0001_1100_1100_0110;     //180pi/512
  assign sin[181]  =  16'b1100_0110_1010_1000;     //181pi/512
  assign cos[181]  =  16'b0001_1100_0110_1100;     //181pi/512
  assign sin[182]  =  16'b1100_0110_0111_1100;     //182pi/512
  assign cos[182]  =  16'b0001_1100_0001_0010;     //182pi/512
  assign sin[183]  =  16'b1100_0110_0101_0000;     //183pi/512
  assign cos[183]  =  16'b0001_1011_1011_0111;     //183pi/512
  assign sin[184]  =  16'b1100_0110_0010_0101;     //184pi/512
  assign cos[184]  =  16'b0001_1011_0101_1101;     //184pi/512
  assign sin[185]  =  16'b1100_0101_1111_1010;     //185pi/512
  assign cos[185]  =  16'b0001_1011_0000_0010;     //185pi/512
  assign sin[186]  =  16'b1100_0101_1101_0000;     //186pi/512
  assign cos[186]  =  16'b0001_1010_1010_0110;     //186pi/512
  assign sin[187]  =  16'b1100_0101_1010_0111;     //187pi/512
  assign cos[187]  =  16'b0001_1010_0100_1011;     //187pi/512
  assign sin[188]  =  16'b1100_0101_0111_1110;     //188pi/512
  assign cos[188]  =  16'b0001_1001_1110_1111;     //188pi/512
  assign sin[189]  =  16'b1100_0101_0101_0101;     //189pi/512
  assign cos[189]  =  16'b0001_1001_1001_0011;     //189pi/512
  assign sin[190]  =  16'b1100_0101_0010_1101;     //190pi/512
  assign cos[190]  =  16'b0001_1001_0011_0111;     //190pi/512
  assign sin[191]  =  16'b1100_0101_0000_0110;     //191pi/512
  assign cos[191]  =  16'b0001_1000_1101_1010;     //191pi/512
  assign sin[192]  =  16'b1100_0100_1101_1111;     //192pi/512
  assign cos[192]  =  16'b0001_1000_0111_1101;     //192pi/512
  assign sin[193]  =  16'b1100_0100_1011_1001;     //193pi/512
  assign cos[193]  =  16'b0001_1000_0010_0000;     //193pi/512
  assign sin[194]  =  16'b1100_0100_1001_0011;     //194pi/512
  assign cos[194]  =  16'b0001_0111_1100_0011;     //194pi/512
  assign sin[195]  =  16'b1100_0100_0110_1110;     //195pi/512
  assign cos[195]  =  16'b0001_0111_0110_0110;     //195pi/512
  assign sin[196]  =  16'b1100_0100_0100_1010;     //196pi/512
  assign cos[196]  =  16'b0001_0111_0000_1000;     //196pi/512
  assign sin[197]  =  16'b1100_0100_0010_0110;     //197pi/512
  assign cos[197]  =  16'b0001_0110_1010_1010;     //197pi/512
  assign sin[198]  =  16'b1100_0100_0000_0011;     //198pi/512
  assign cos[198]  =  16'b0001_0110_0100_1100;     //198pi/512
  assign sin[199]  =  16'b1100_0011_1110_0000;     //199pi/512
  assign cos[199]  =  16'b0001_0101_1110_1110;     //199pi/512
  assign sin[200]  =  16'b1100_0011_1011_1110;     //200pi/512
  assign cos[200]  =  16'b0001_0101_1000_1111;     //200pi/512
  assign sin[201]  =  16'b1100_0011_1001_1100;     //201pi/512
  assign cos[201]  =  16'b0001_0101_0011_0000;     //201pi/512
  assign sin[202]  =  16'b1100_0011_0111_1011;     //202pi/512
  assign cos[202]  =  16'b0001_0100_1101_0001;     //202pi/512
  assign sin[203]  =  16'b1100_0011_0101_1011;     //203pi/512
  assign cos[203]  =  16'b0001_0100_0111_0010;     //203pi/512
  assign sin[204]  =  16'b1100_0011_0011_1011;     //204pi/512
  assign cos[204]  =  16'b0001_0100_0001_0011;     //204pi/512
  assign sin[205]  =  16'b1100_0011_0001_1100;     //205pi/512
  assign cos[205]  =  16'b0001_0011_1011_0011;     //205pi/512
  assign sin[206]  =  16'b1100_0010_1111_1101;     //206pi/512
  assign cos[206]  =  16'b0001_0011_0101_0100;     //206pi/512
  assign sin[207]  =  16'b1100_0010_1101_1111;     //207pi/512
  assign cos[207]  =  16'b0001_0010_1111_0100;     //207pi/512
  assign sin[208]  =  16'b1100_0010_1100_0001;     //208pi/512
  assign cos[208]  =  16'b0001_0010_1001_0100;     //208pi/512
  assign sin[209]  =  16'b1100_0010_1010_0101;     //209pi/512
  assign cos[209]  =  16'b0001_0010_0011_0011;     //209pi/512
  assign sin[210]  =  16'b1100_0010_1000_1000;     //210pi/512
  assign cos[210]  =  16'b0001_0001_1101_0011;     //210pi/512
  assign sin[211]  =  16'b1100_0010_0110_1101;     //211pi/512
  assign cos[211]  =  16'b0001_0001_0111_0010;     //211pi/512
  assign sin[212]  =  16'b1100_0010_0101_0001;     //212pi/512
  assign cos[212]  =  16'b0001_0001_0001_0001;     //212pi/512
  assign sin[213]  =  16'b1100_0010_0011_0111;     //213pi/512
  assign cos[213]  =  16'b0001_0000_1011_0000;     //213pi/512
  assign sin[214]  =  16'b1100_0010_0001_1101;     //214pi/512
  assign cos[214]  =  16'b0001_0000_0100_1111;     //214pi/512
  assign sin[215]  =  16'b1100_0010_0000_0100;     //215pi/512
  assign cos[215]  =  16'b0000_1111_1110_1110;     //215pi/512
  assign sin[216]  =  16'b1100_0001_1110_1011;     //216pi/512
  assign cos[216]  =  16'b0000_1111_1000_1100;     //216pi/512
  assign sin[217]  =  16'b1100_0001_1101_0011;     //217pi/512
  assign cos[217]  =  16'b0000_1111_0010_1011;     //217pi/512
  assign sin[218]  =  16'b1100_0001_1011_1011;     //218pi/512
  assign cos[218]  =  16'b0000_1110_1100_1001;     //218pi/512
  assign sin[219]  =  16'b1100_0001_1010_0100;     //219pi/512
  assign cos[219]  =  16'b0000_1110_0110_0111;     //219pi/512
  assign sin[220]  =  16'b1100_0001_1000_1110;     //220pi/512
  assign cos[220]  =  16'b0000_1110_0000_0101;     //220pi/512
  assign sin[221]  =  16'b1100_0001_0111_1000;     //221pi/512
  assign cos[221]  =  16'b0000_1101_1010_0011;     //221pi/512
  assign sin[222]  =  16'b1100_0001_0110_0011;     //222pi/512
  assign cos[222]  =  16'b0000_1101_0100_0001;     //222pi/512
  assign sin[223]  =  16'b1100_0001_0100_1111;     //223pi/512
  assign cos[223]  =  16'b0000_1100_1101_1110;     //223pi/512
  assign sin[224]  =  16'b1100_0001_0011_1011;     //224pi/512
  assign cos[224]  =  16'b0000_1100_0111_1100;     //224pi/512
  assign sin[225]  =  16'b1100_0001_0010_1000;     //225pi/512
  assign cos[225]  =  16'b0000_1100_0001_1001;     //225pi/512
  assign sin[226]  =  16'b1100_0001_0001_0101;     //226pi/512
  assign cos[226]  =  16'b0000_1011_1011_0110;     //226pi/512
  assign sin[227]  =  16'b1100_0001_0000_0011;     //227pi/512
  assign cos[227]  =  16'b0000_1011_0101_0100;     //227pi/512
  assign sin[228]  =  16'b1100_0000_1111_0001;     //228pi/512
  assign cos[228]  =  16'b0000_1010_1111_0001;     //228pi/512
  assign sin[229]  =  16'b1100_0000_1110_0000;     //229pi/512
  assign cos[229]  =  16'b0000_1010_1000_1101;     //229pi/512
  assign sin[230]  =  16'b1100_0000_1101_0000;     //230pi/512
  assign cos[230]  =  16'b0000_1010_0010_1010;     //230pi/512
  assign sin[231]  =  16'b1100_0000_1100_0000;     //231pi/512
  assign cos[231]  =  16'b0000_1001_1100_0111;     //231pi/512
  assign sin[232]  =  16'b1100_0000_1011_0001;     //232pi/512
  assign cos[232]  =  16'b0000_1001_0110_0100;     //232pi/512
  assign sin[233]  =  16'b1100_0000_1010_0011;     //233pi/512
  assign cos[233]  =  16'b0000_1001_0000_0000;     //233pi/512
  assign sin[234]  =  16'b1100_0000_1001_0101;     //234pi/512
  assign cos[234]  =  16'b0000_1000_1001_1100;     //234pi/512
  assign sin[235]  =  16'b1100_0000_1000_1000;     //235pi/512
  assign cos[235]  =  16'b0000_1000_0011_1001;     //235pi/512
  assign sin[236]  =  16'b1100_0000_0111_1011;     //236pi/512
  assign cos[236]  =  16'b0000_0111_1101_0101;     //236pi/512
  assign sin[237]  =  16'b1100_0000_0110_1111;     //237pi/512
  assign cos[237]  =  16'b0000_0111_0111_0001;     //237pi/512
  assign sin[238]  =  16'b1100_0000_0110_0100;     //238pi/512
  assign cos[238]  =  16'b0000_0111_0000_1101;     //238pi/512
  assign sin[239]  =  16'b1100_0000_0101_1001;     //239pi/512
  assign cos[239]  =  16'b0000_0110_1010_1001;     //239pi/512
  assign sin[240]  =  16'b1100_0000_0100_1111;     //240pi/512
  assign cos[240]  =  16'b0000_0110_0100_0101;     //240pi/512
  assign sin[241]  =  16'b1100_0000_0100_0101;     //241pi/512
  assign cos[241]  =  16'b0000_0101_1110_0001;     //241pi/512
  assign sin[242]  =  16'b1100_0000_0011_1100;     //242pi/512
  assign cos[242]  =  16'b0000_0101_0111_1101;     //242pi/512
  assign sin[243]  =  16'b1100_0000_0011_0100;     //243pi/512
  assign cos[243]  =  16'b0000_0101_0001_1001;     //243pi/512
  assign sin[244]  =  16'b1100_0000_0010_1100;     //244pi/512
  assign cos[244]  =  16'b0000_0100_1011_0101;     //244pi/512
  assign sin[245]  =  16'b1100_0000_0010_0101;     //245pi/512
  assign cos[245]  =  16'b0000_0100_0101_0001;     //245pi/512
  assign sin[246]  =  16'b1100_0000_0001_1111;     //246pi/512
  assign cos[246]  =  16'b0000_0011_1110_1100;     //246pi/512
  assign sin[247]  =  16'b1100_0000_0001_1001;     //247pi/512
  assign cos[247]  =  16'b0000_0011_1000_1000;     //247pi/512
  assign sin[248]  =  16'b1100_0000_0001_0100;     //248pi/512
  assign cos[248]  =  16'b0000_0011_0010_0011;     //248pi/512
  assign sin[249]  =  16'b1100_0000_0000_1111;     //249pi/512
  assign cos[249]  =  16'b0000_0010_1011_1111;     //249pi/512
  assign sin[250]  =  16'b1100_0000_0000_1011;     //250pi/512
  assign cos[250]  =  16'b0000_0010_0101_1011;     //250pi/512
  assign sin[251]  =  16'b1100_0000_0000_1000;     //251pi/512
  assign cos[251]  =  16'b0000_0001_1111_0110;     //251pi/512
  assign sin[252]  =  16'b1100_0000_0000_0101;     //252pi/512
  assign cos[252]  =  16'b0000_0001_1001_0010;     //252pi/512
  assign sin[253]  =  16'b1100_0000_0000_0011;     //253pi/512
  assign cos[253]  =  16'b0000_0001_0010_1101;     //253pi/512
  assign sin[254]  =  16'b1100_0000_0000_0001;     //254pi/512
  assign cos[254]  =  16'b0000_0000_1100_1001;     //254pi/512
  assign sin[255]  =  16'b1100_0000_0000_0000;     //255pi/512
  assign cos[255]  =  16'b0000_0000_0110_0100;     //255pi/512
  assign sin[256]  =  16'b1100_0000_0000_0000;     //256pi/512
  assign cos[256]  =  16'b0000_0000_0000_0000;     //256pi/512
  assign sin[257]  =  16'b1100_0000_0000_0000;     //257pi/512
  assign cos[257]  =  16'b1111_1111_1001_1011;     //257pi/512
  assign sin[258]  =  16'b1100_0000_0000_0001;     //258pi/512
  assign cos[258]  =  16'b1111_1111_0011_0111;     //258pi/512
  assign sin[259]  =  16'b1100_0000_0000_0011;     //259pi/512
  assign cos[259]  =  16'b1111_1110_1101_0010;     //259pi/512
  assign sin[260]  =  16'b1100_0000_0000_0101;     //260pi/512
  assign cos[260]  =  16'b1111_1110_0110_1110;     //260pi/512
  assign sin[261]  =  16'b1100_0000_0000_1000;     //261pi/512
  assign cos[261]  =  16'b1111_1110_0000_1001;     //261pi/512
  assign sin[262]  =  16'b1100_0000_0000_1011;     //262pi/512
  assign cos[262]  =  16'b1111_1101_1010_0101;     //262pi/512
  assign sin[263]  =  16'b1100_0000_0000_1111;     //263pi/512
  assign cos[263]  =  16'b1111_1101_0100_0000;     //263pi/512
  assign sin[264]  =  16'b1100_0000_0001_0100;     //264pi/512
  assign cos[264]  =  16'b1111_1100_1101_1100;     //264pi/512
  assign sin[265]  =  16'b1100_0000_0001_1001;     //265pi/512
  assign cos[265]  =  16'b1111_1100_0111_1000;     //265pi/512
  assign sin[266]  =  16'b1100_0000_0001_1111;     //266pi/512
  assign cos[266]  =  16'b1111_1100_0001_0011;     //266pi/512
  assign sin[267]  =  16'b1100_0000_0010_0101;     //267pi/512
  assign cos[267]  =  16'b1111_1011_1010_1111;     //267pi/512
  assign sin[268]  =  16'b1100_0000_0010_1100;     //268pi/512
  assign cos[268]  =  16'b1111_1011_0100_1011;     //268pi/512
  assign sin[269]  =  16'b1100_0000_0011_0100;     //269pi/512
  assign cos[269]  =  16'b1111_1010_1110_0110;     //269pi/512
  assign sin[270]  =  16'b1100_0000_0011_1100;     //270pi/512
  assign cos[270]  =  16'b1111_1010_1000_0010;     //270pi/512
  assign sin[271]  =  16'b1100_0000_0100_0101;     //271pi/512
  assign cos[271]  =  16'b1111_1010_0001_1110;     //271pi/512
  assign sin[272]  =  16'b1100_0000_0100_1111;     //272pi/512
  assign cos[272]  =  16'b1111_1001_1011_1010;     //272pi/512
  assign sin[273]  =  16'b1100_0000_0101_1001;     //273pi/512
  assign cos[273]  =  16'b1111_1001_0101_0110;     //273pi/512
  assign sin[274]  =  16'b1100_0000_0110_0100;     //274pi/512
  assign cos[274]  =  16'b1111_1000_1111_0010;     //274pi/512
  assign sin[275]  =  16'b1100_0000_0110_1111;     //275pi/512
  assign cos[275]  =  16'b1111_1000_1000_1110;     //275pi/512
  assign sin[276]  =  16'b1100_0000_0111_1011;     //276pi/512
  assign cos[276]  =  16'b1111_1000_0010_1010;     //276pi/512
  assign sin[277]  =  16'b1100_0000_1000_1000;     //277pi/512
  assign cos[277]  =  16'b1111_0111_1100_0111;     //277pi/512
  assign sin[278]  =  16'b1100_0000_1001_0101;     //278pi/512
  assign cos[278]  =  16'b1111_0111_0110_0011;     //278pi/512
  assign sin[279]  =  16'b1100_0000_1010_0011;     //279pi/512
  assign cos[279]  =  16'b1111_0110_1111_1111;     //279pi/512
  assign sin[280]  =  16'b1100_0000_1011_0001;     //280pi/512
  assign cos[280]  =  16'b1111_0110_1001_1100;     //280pi/512
  assign sin[281]  =  16'b1100_0000_1100_0000;     //281pi/512
  assign cos[281]  =  16'b1111_0110_0011_1001;     //281pi/512
  assign sin[282]  =  16'b1100_0000_1101_0000;     //282pi/512
  assign cos[282]  =  16'b1111_0101_1101_0101;     //282pi/512
  assign sin[283]  =  16'b1100_0000_1110_0000;     //283pi/512
  assign cos[283]  =  16'b1111_0101_0111_0010;     //283pi/512
  assign sin[284]  =  16'b1100_0000_1111_0001;     //284pi/512
  assign cos[284]  =  16'b1111_0101_0000_1111;     //284pi/512
  assign sin[285]  =  16'b1100_0001_0000_0011;     //285pi/512
  assign cos[285]  =  16'b1111_0100_1010_1100;     //285pi/512
  assign sin[286]  =  16'b1100_0001_0001_0101;     //286pi/512
  assign cos[286]  =  16'b1111_0100_0100_1001;     //286pi/512
  assign sin[287]  =  16'b1100_0001_0010_1000;     //287pi/512
  assign cos[287]  =  16'b1111_0011_1110_0110;     //287pi/512
  assign sin[288]  =  16'b1100_0001_0011_1011;     //288pi/512
  assign cos[288]  =  16'b1111_0011_1000_0100;     //288pi/512
  assign sin[289]  =  16'b1100_0001_0100_1111;     //289pi/512
  assign cos[289]  =  16'b1111_0011_0010_0001;     //289pi/512
  assign sin[290]  =  16'b1100_0001_0110_0011;     //290pi/512
  assign cos[290]  =  16'b1111_0010_1011_1111;     //290pi/512
  assign sin[291]  =  16'b1100_0001_0111_1000;     //291pi/512
  assign cos[291]  =  16'b1111_0010_0101_1100;     //291pi/512
  assign sin[292]  =  16'b1100_0001_1000_1110;     //292pi/512
  assign cos[292]  =  16'b1111_0001_1111_1010;     //292pi/512
  assign sin[293]  =  16'b1100_0001_1010_0100;     //293pi/512
  assign cos[293]  =  16'b1111_0001_1001_1000;     //293pi/512
  assign sin[294]  =  16'b1100_0001_1011_1011;     //294pi/512
  assign cos[294]  =  16'b1111_0001_0011_0110;     //294pi/512
  assign sin[295]  =  16'b1100_0001_1101_0011;     //295pi/512
  assign cos[295]  =  16'b1111_0000_1101_0101;     //295pi/512
  assign sin[296]  =  16'b1100_0001_1110_1011;     //296pi/512
  assign cos[296]  =  16'b1111_0000_0111_0011;     //296pi/512
  assign sin[297]  =  16'b1100_0010_0000_0100;     //297pi/512
  assign cos[297]  =  16'b1111_0000_0001_0010;     //297pi/512
  assign sin[298]  =  16'b1100_0010_0001_1101;     //298pi/512
  assign cos[298]  =  16'b1110_1111_1011_0000;     //298pi/512
  assign sin[299]  =  16'b1100_0010_0011_0111;     //299pi/512
  assign cos[299]  =  16'b1110_1111_0100_1111;     //299pi/512
  assign sin[300]  =  16'b1100_0010_0101_0001;     //300pi/512
  assign cos[300]  =  16'b1110_1110_1110_1110;     //300pi/512
  assign sin[301]  =  16'b1100_0010_0110_1101;     //301pi/512
  assign cos[301]  =  16'b1110_1110_1000_1101;     //301pi/512
  assign sin[302]  =  16'b1100_0010_1000_1000;     //302pi/512
  assign cos[302]  =  16'b1110_1110_0010_1101;     //302pi/512
  assign sin[303]  =  16'b1100_0010_1010_0101;     //303pi/512
  assign cos[303]  =  16'b1110_1101_1100_1100;     //303pi/512
  assign sin[304]  =  16'b1100_0010_1100_0001;     //304pi/512
  assign cos[304]  =  16'b1110_1101_0110_1100;     //304pi/512
  assign sin[305]  =  16'b1100_0010_1101_1111;     //305pi/512
  assign cos[305]  =  16'b1110_1101_0000_1100;     //305pi/512
  assign sin[306]  =  16'b1100_0010_1111_1101;     //306pi/512
  assign cos[306]  =  16'b1110_1100_1010_1100;     //306pi/512
  assign sin[307]  =  16'b1100_0011_0001_1100;     //307pi/512
  assign cos[307]  =  16'b1110_1100_0100_1100;     //307pi/512
  assign sin[308]  =  16'b1100_0011_0011_1011;     //308pi/512
  assign cos[308]  =  16'b1110_1011_1110_1101;     //308pi/512
  assign sin[309]  =  16'b1100_0011_0101_1011;     //309pi/512
  assign cos[309]  =  16'b1110_1011_1000_1101;     //309pi/512
  assign sin[310]  =  16'b1100_0011_0111_1011;     //310pi/512
  assign cos[310]  =  16'b1110_1011_0010_1110;     //310pi/512
  assign sin[311]  =  16'b1100_0011_1001_1100;     //311pi/512
  assign cos[311]  =  16'b1110_1010_1100_1111;     //311pi/512
  assign sin[312]  =  16'b1100_0011_1011_1110;     //312pi/512
  assign cos[312]  =  16'b1110_1010_0111_0000;     //312pi/512
  assign sin[313]  =  16'b1100_0011_1110_0000;     //313pi/512
  assign cos[313]  =  16'b1110_1010_0001_0010;     //313pi/512
  assign sin[314]  =  16'b1100_0100_0000_0011;     //314pi/512
  assign cos[314]  =  16'b1110_1001_1011_0100;     //314pi/512
  assign sin[315]  =  16'b1100_0100_0010_0110;     //315pi/512
  assign cos[315]  =  16'b1110_1001_0101_0101;     //315pi/512
  assign sin[316]  =  16'b1100_0100_0100_1010;     //316pi/512
  assign cos[316]  =  16'b1110_1000_1111_0111;     //316pi/512
  assign sin[317]  =  16'b1100_0100_0110_1110;     //317pi/512
  assign cos[317]  =  16'b1110_1000_1001_1010;     //317pi/512
  assign sin[318]  =  16'b1100_0100_1001_0011;     //318pi/512
  assign cos[318]  =  16'b1110_1000_0011_1100;     //318pi/512
  assign sin[319]  =  16'b1100_0100_1011_1001;     //319pi/512
  assign cos[319]  =  16'b1110_0111_1101_1111;     //319pi/512
  assign sin[320]  =  16'b1100_0100_1101_1111;     //320pi/512
  assign cos[320]  =  16'b1110_0111_1000_0010;     //320pi/512
  assign sin[321]  =  16'b1100_0101_0000_0110;     //321pi/512
  assign cos[321]  =  16'b1110_0111_0010_0101;     //321pi/512
  assign sin[322]  =  16'b1100_0101_0010_1101;     //322pi/512
  assign cos[322]  =  16'b1110_0110_1100_1001;     //322pi/512
  assign sin[323]  =  16'b1100_0101_0101_0101;     //323pi/512
  assign cos[323]  =  16'b1110_0110_0110_1101;     //323pi/512
  assign sin[324]  =  16'b1100_0101_0111_1110;     //324pi/512
  assign cos[324]  =  16'b1110_0110_0001_0001;     //324pi/512
  assign sin[325]  =  16'b1100_0101_1010_0111;     //325pi/512
  assign cos[325]  =  16'b1110_0101_1011_0101;     //325pi/512
  assign sin[326]  =  16'b1100_0101_1101_0000;     //326pi/512
  assign cos[326]  =  16'b1110_0101_0101_1001;     //326pi/512
  assign sin[327]  =  16'b1100_0101_1111_1010;     //327pi/512
  assign cos[327]  =  16'b1110_0100_1111_1110;     //327pi/512
  assign sin[328]  =  16'b1100_0110_0010_0101;     //328pi/512
  assign cos[328]  =  16'b1110_0100_1010_0011;     //328pi/512
  assign sin[329]  =  16'b1100_0110_0101_0000;     //329pi/512
  assign cos[329]  =  16'b1110_0100_0100_1000;     //329pi/512
  assign sin[330]  =  16'b1100_0110_0111_1100;     //330pi/512
  assign cos[330]  =  16'b1110_0011_1110_1110;     //330pi/512
  assign sin[331]  =  16'b1100_0110_1010_1000;     //331pi/512
  assign cos[331]  =  16'b1110_0011_1001_0100;     //331pi/512
  assign sin[332]  =  16'b1100_0110_1101_0101;     //332pi/512
  assign cos[332]  =  16'b1110_0011_0011_1010;     //332pi/512
  assign sin[333]  =  16'b1100_0111_0000_0011;     //333pi/512
  assign cos[333]  =  16'b1110_0010_1110_0000;     //333pi/512
  assign sin[334]  =  16'b1100_0111_0011_0001;     //334pi/512
  assign cos[334]  =  16'b1110_0010_1000_0111;     //334pi/512
  assign sin[335]  =  16'b1100_0111_0101_1111;     //335pi/512
  assign cos[335]  =  16'b1110_0010_0010_1101;     //335pi/512
  assign sin[336]  =  16'b1100_0111_1000_1111;     //336pi/512
  assign cos[336]  =  16'b1110_0001_1101_0101;     //336pi/512
  assign sin[337]  =  16'b1100_0111_1011_1110;     //337pi/512
  assign cos[337]  =  16'b1110_0001_0111_1100;     //337pi/512
  assign sin[338]  =  16'b1100_0111_1110_1110;     //338pi/512
  assign cos[338]  =  16'b1110_0001_0010_0100;     //338pi/512
  assign sin[339]  =  16'b1100_1000_0001_1111;     //339pi/512
  assign cos[339]  =  16'b1110_0000_1100_1100;     //339pi/512
  assign sin[340]  =  16'b1100_1000_0101_0000;     //340pi/512
  assign cos[340]  =  16'b1110_0000_0111_0100;     //340pi/512
  assign sin[341]  =  16'b1100_1000_1000_0010;     //341pi/512
  assign cos[341]  =  16'b1110_0000_0001_1101;     //341pi/512
  assign sin[342]  =  16'b1100_1000_1011_0101;     //342pi/512
  assign cos[342]  =  16'b1101_1111_1100_0110;     //342pi/512
  assign sin[343]  =  16'b1100_1000_1110_1000;     //343pi/512
  assign cos[343]  =  16'b1101_1111_0110_1111;     //343pi/512
  assign sin[344]  =  16'b1100_1001_0001_1011;     //344pi/512
  assign cos[344]  =  16'b1101_1111_0001_1001;     //344pi/512
  assign sin[345]  =  16'b1100_1001_0100_1111;     //345pi/512
  assign cos[345]  =  16'b1101_1110_1100_0011;     //345pi/512
  assign sin[346]  =  16'b1100_1001_1000_0011;     //346pi/512
  assign cos[346]  =  16'b1101_1110_0110_1101;     //346pi/512
  assign sin[347]  =  16'b1100_1001_1011_1000;     //347pi/512
  assign cos[347]  =  16'b1101_1110_0001_1000;     //347pi/512
  assign sin[348]  =  16'b1100_1001_1110_1110;     //348pi/512
  assign cos[348]  =  16'b1101_1101_1100_0011;     //348pi/512
  assign sin[349]  =  16'b1100_1010_0010_0100;     //349pi/512
  assign cos[349]  =  16'b1101_1101_0110_1110;     //349pi/512
  assign sin[350]  =  16'b1100_1010_0101_1011;     //350pi/512
  assign cos[350]  =  16'b1101_1101_0001_1001;     //350pi/512
  assign sin[351]  =  16'b1100_1010_1001_0010;     //351pi/512
  assign cos[351]  =  16'b1101_1100_1100_0101;     //351pi/512
  assign sin[352]  =  16'b1100_1010_1100_1001;     //352pi/512
  assign cos[352]  =  16'b1101_1100_0111_0010;     //352pi/512
  assign sin[353]  =  16'b1100_1011_0000_0001;     //353pi/512
  assign cos[353]  =  16'b1101_1100_0001_1110;     //353pi/512
  assign sin[354]  =  16'b1100_1011_0011_1010;     //354pi/512
  assign cos[354]  =  16'b1101_1011_1100_1011;     //354pi/512
  assign sin[355]  =  16'b1100_1011_0111_0011;     //355pi/512
  assign cos[355]  =  16'b1101_1011_0111_1000;     //355pi/512
  assign sin[356]  =  16'b1100_1011_1010_1101;     //356pi/512
  assign cos[356]  =  16'b1101_1011_0010_0110;     //356pi/512
  assign sin[357]  =  16'b1100_1011_1110_0111;     //357pi/512
  assign cos[357]  =  16'b1101_1010_1101_0100;     //357pi/512
  assign sin[358]  =  16'b1100_1100_0010_0001;     //358pi/512
  assign cos[358]  =  16'b1101_1010_1000_0010;     //358pi/512
  assign sin[359]  =  16'b1100_1100_0101_1101;     //359pi/512
  assign cos[359]  =  16'b1101_1010_0011_0001;     //359pi/512
  assign sin[360]  =  16'b1100_1100_1001_1000;     //360pi/512
  assign cos[360]  =  16'b1101_1001_1110_0000;     //360pi/512
  assign sin[361]  =  16'b1100_1100_1101_0100;     //361pi/512
  assign cos[361]  =  16'b1101_1001_1000_1111;     //361pi/512
  assign sin[362]  =  16'b1100_1101_0001_0001;     //362pi/512
  assign cos[362]  =  16'b1101_1001_0011_1111;     //362pi/512
  assign sin[363]  =  16'b1100_1101_0100_1110;     //363pi/512
  assign cos[363]  =  16'b1101_1000_1110_1111;     //363pi/512
  assign sin[364]  =  16'b1100_1101_1000_1100;     //364pi/512
  assign cos[364]  =  16'b1101_1000_1010_0000;     //364pi/512
  assign sin[365]  =  16'b1100_1101_1100_1010;     //365pi/512
  assign cos[365]  =  16'b1101_1000_0101_0001;     //365pi/512
  assign sin[366]  =  16'b1100_1110_0000_1000;     //366pi/512
  assign cos[366]  =  16'b1101_1000_0000_0010;     //366pi/512
  assign sin[367]  =  16'b1100_1110_0100_0111;     //367pi/512
  assign cos[367]  =  16'b1101_0111_1011_0100;     //367pi/512
  assign sin[368]  =  16'b1100_1110_1000_0111;     //368pi/512
  assign cos[368]  =  16'b1101_0111_0110_0110;     //368pi/512
  assign sin[369]  =  16'b1100_1110_1100_0111;     //369pi/512
  assign cos[369]  =  16'b1101_0111_0001_1001;     //369pi/512
  assign sin[370]  =  16'b1100_1111_0000_0111;     //370pi/512
  assign cos[370]  =  16'b1101_0110_1100_1011;     //370pi/512
  assign sin[371]  =  16'b1100_1111_0100_1000;     //371pi/512
  assign cos[371]  =  16'b1101_0110_0111_1111;     //371pi/512
  assign sin[372]  =  16'b1100_1111_1000_1010;     //372pi/512
  assign cos[372]  =  16'b1101_0110_0011_0010;     //372pi/512
  assign sin[373]  =  16'b1100_1111_1100_1100;     //373pi/512
  assign cos[373]  =  16'b1101_0101_1110_0110;     //373pi/512
  assign sin[374]  =  16'b1101_0000_0000_1110;     //374pi/512
  assign cos[374]  =  16'b1101_0101_1001_1011;     //374pi/512
  assign sin[375]  =  16'b1101_0000_0101_0001;     //375pi/512
  assign cos[375]  =  16'b1101_0101_0101_0000;     //375pi/512
  assign sin[376]  =  16'b1101_0000_1001_0100;     //376pi/512
  assign cos[376]  =  16'b1101_0101_0000_0101;     //376pi/512
  assign sin[377]  =  16'b1101_0000_1101_1000;     //377pi/512
  assign cos[377]  =  16'b1101_0100_1011_1011;     //377pi/512
  assign sin[378]  =  16'b1101_0001_0001_1100;     //378pi/512
  assign cos[378]  =  16'b1101_0100_0111_0001;     //378pi/512
  assign sin[379]  =  16'b1101_0001_0110_0001;     //379pi/512
  assign cos[379]  =  16'b1101_0100_0010_1000;     //379pi/512
  assign sin[380]  =  16'b1101_0001_1010_0110;     //380pi/512
  assign cos[380]  =  16'b1101_0011_1101_1111;     //380pi/512
  assign sin[381]  =  16'b1101_0001_1110_1011;     //381pi/512
  assign cos[381]  =  16'b1101_0011_1001_0110;     //381pi/512
  assign sin[382]  =  16'b1101_0010_0011_0001;     //382pi/512
  assign cos[382]  =  16'b1101_0011_0100_1110;     //382pi/512
  assign sin[383]  =  16'b1101_0010_0111_1000;     //383pi/512
  assign cos[383]  =  16'b1101_0011_0000_0110;     //383pi/512
  assign sin[384]  =  16'b1101_0010_1011_1111;     //384pi/512
  assign cos[384]  =  16'b1101_0010_1011_1111;     //384pi/512
  assign sin[385]  =  16'b1101_0011_0000_0110;     //385pi/512
  assign cos[385]  =  16'b1101_0010_0111_1000;     //385pi/512
  assign sin[386]  =  16'b1101_0011_0100_1110;     //386pi/512
  assign cos[386]  =  16'b1101_0010_0011_0001;     //386pi/512
  assign sin[387]  =  16'b1101_0011_1001_0110;     //387pi/512
  assign cos[387]  =  16'b1101_0001_1110_1011;     //387pi/512
  assign sin[388]  =  16'b1101_0011_1101_1111;     //388pi/512
  assign cos[388]  =  16'b1101_0001_1010_0110;     //388pi/512
  assign sin[389]  =  16'b1101_0100_0010_1000;     //389pi/512
  assign cos[389]  =  16'b1101_0001_0110_0001;     //389pi/512
  assign sin[390]  =  16'b1101_0100_0111_0001;     //390pi/512
  assign cos[390]  =  16'b1101_0001_0001_1100;     //390pi/512
  assign sin[391]  =  16'b1101_0100_1011_1011;     //391pi/512
  assign cos[391]  =  16'b1101_0000_1101_1000;     //391pi/512
  assign sin[392]  =  16'b1101_0101_0000_0101;     //392pi/512
  assign cos[392]  =  16'b1101_0000_1001_0100;     //392pi/512
  assign sin[393]  =  16'b1101_0101_0101_0000;     //393pi/512
  assign cos[393]  =  16'b1101_0000_0101_0001;     //393pi/512
  assign sin[394]  =  16'b1101_0101_1001_1011;     //394pi/512
  assign cos[394]  =  16'b1101_0000_0000_1110;     //394pi/512
  assign sin[395]  =  16'b1101_0101_1110_0110;     //395pi/512
  assign cos[395]  =  16'b1100_1111_1100_1100;     //395pi/512
  assign sin[396]  =  16'b1101_0110_0011_0010;     //396pi/512
  assign cos[396]  =  16'b1100_1111_1000_1010;     //396pi/512
  assign sin[397]  =  16'b1101_0110_0111_1111;     //397pi/512
  assign cos[397]  =  16'b1100_1111_0100_1000;     //397pi/512
  assign sin[398]  =  16'b1101_0110_1100_1011;     //398pi/512
  assign cos[398]  =  16'b1100_1111_0000_0111;     //398pi/512
  assign sin[399]  =  16'b1101_0111_0001_1001;     //399pi/512
  assign cos[399]  =  16'b1100_1110_1100_0111;     //399pi/512
  assign sin[400]  =  16'b1101_0111_0110_0110;     //400pi/512
  assign cos[400]  =  16'b1100_1110_1000_0111;     //400pi/512
  assign sin[401]  =  16'b1101_0111_1011_0100;     //401pi/512
  assign cos[401]  =  16'b1100_1110_0100_0111;     //401pi/512
  assign sin[402]  =  16'b1101_1000_0000_0010;     //402pi/512
  assign cos[402]  =  16'b1100_1110_0000_1000;     //402pi/512
  assign sin[403]  =  16'b1101_1000_0101_0001;     //403pi/512
  assign cos[403]  =  16'b1100_1101_1100_1010;     //403pi/512
  assign sin[404]  =  16'b1101_1000_1010_0000;     //404pi/512
  assign cos[404]  =  16'b1100_1101_1000_1100;     //404pi/512
  assign sin[405]  =  16'b1101_1000_1110_1111;     //405pi/512
  assign cos[405]  =  16'b1100_1101_0100_1110;     //405pi/512
  assign sin[406]  =  16'b1101_1001_0011_1111;     //406pi/512
  assign cos[406]  =  16'b1100_1101_0001_0001;     //406pi/512
  assign sin[407]  =  16'b1101_1001_1000_1111;     //407pi/512
  assign cos[407]  =  16'b1100_1100_1101_0100;     //407pi/512
  assign sin[408]  =  16'b1101_1001_1110_0000;     //408pi/512
  assign cos[408]  =  16'b1100_1100_1001_1000;     //408pi/512
  assign sin[409]  =  16'b1101_1010_0011_0001;     //409pi/512
  assign cos[409]  =  16'b1100_1100_0101_1101;     //409pi/512
  assign sin[410]  =  16'b1101_1010_1000_0010;     //410pi/512
  assign cos[410]  =  16'b1100_1100_0010_0001;     //410pi/512
  assign sin[411]  =  16'b1101_1010_1101_0100;     //411pi/512
  assign cos[411]  =  16'b1100_1011_1110_0111;     //411pi/512
  assign sin[412]  =  16'b1101_1011_0010_0110;     //412pi/512
  assign cos[412]  =  16'b1100_1011_1010_1101;     //412pi/512
  assign sin[413]  =  16'b1101_1011_0111_1000;     //413pi/512
  assign cos[413]  =  16'b1100_1011_0111_0011;     //413pi/512
  assign sin[414]  =  16'b1101_1011_1100_1011;     //414pi/512
  assign cos[414]  =  16'b1100_1011_0011_1010;     //414pi/512
  assign sin[415]  =  16'b1101_1100_0001_1110;     //415pi/512
  assign cos[415]  =  16'b1100_1011_0000_0001;     //415pi/512
  assign sin[416]  =  16'b1101_1100_0111_0010;     //416pi/512
  assign cos[416]  =  16'b1100_1010_1100_1001;     //416pi/512
  assign sin[417]  =  16'b1101_1100_1100_0101;     //417pi/512
  assign cos[417]  =  16'b1100_1010_1001_0010;     //417pi/512
  assign sin[418]  =  16'b1101_1101_0001_1001;     //418pi/512
  assign cos[418]  =  16'b1100_1010_0101_1011;     //418pi/512
  assign sin[419]  =  16'b1101_1101_0110_1110;     //419pi/512
  assign cos[419]  =  16'b1100_1010_0010_0100;     //419pi/512
  assign sin[420]  =  16'b1101_1101_1100_0011;     //420pi/512
  assign cos[420]  =  16'b1100_1001_1110_1110;     //420pi/512
  assign sin[421]  =  16'b1101_1110_0001_1000;     //421pi/512
  assign cos[421]  =  16'b1100_1001_1011_1000;     //421pi/512
  assign sin[422]  =  16'b1101_1110_0110_1101;     //422pi/512
  assign cos[422]  =  16'b1100_1001_1000_0011;     //422pi/512
  assign sin[423]  =  16'b1101_1110_1100_0011;     //423pi/512
  assign cos[423]  =  16'b1100_1001_0100_1111;     //423pi/512
  assign sin[424]  =  16'b1101_1111_0001_1001;     //424pi/512
  assign cos[424]  =  16'b1100_1001_0001_1011;     //424pi/512
  assign sin[425]  =  16'b1101_1111_0110_1111;     //425pi/512
  assign cos[425]  =  16'b1100_1000_1110_1000;     //425pi/512
  assign sin[426]  =  16'b1101_1111_1100_0110;     //426pi/512
  assign cos[426]  =  16'b1100_1000_1011_0101;     //426pi/512
  assign sin[427]  =  16'b1110_0000_0001_1101;     //427pi/512
  assign cos[427]  =  16'b1100_1000_1000_0010;     //427pi/512
  assign sin[428]  =  16'b1110_0000_0111_0100;     //428pi/512
  assign cos[428]  =  16'b1100_1000_0101_0000;     //428pi/512
  assign sin[429]  =  16'b1110_0000_1100_1100;     //429pi/512
  assign cos[429]  =  16'b1100_1000_0001_1111;     //429pi/512
  assign sin[430]  =  16'b1110_0001_0010_0100;     //430pi/512
  assign cos[430]  =  16'b1100_0111_1110_1110;     //430pi/512
  assign sin[431]  =  16'b1110_0001_0111_1100;     //431pi/512
  assign cos[431]  =  16'b1100_0111_1011_1110;     //431pi/512
  assign sin[432]  =  16'b1110_0001_1101_0101;     //432pi/512
  assign cos[432]  =  16'b1100_0111_1000_1111;     //432pi/512
  assign sin[433]  =  16'b1110_0010_0010_1101;     //433pi/512
  assign cos[433]  =  16'b1100_0111_0101_1111;     //433pi/512
  assign sin[434]  =  16'b1110_0010_1000_0111;     //434pi/512
  assign cos[434]  =  16'b1100_0111_0011_0001;     //434pi/512
  assign sin[435]  =  16'b1110_0010_1110_0000;     //435pi/512
  assign cos[435]  =  16'b1100_0111_0000_0011;     //435pi/512
  assign sin[436]  =  16'b1110_0011_0011_1010;     //436pi/512
  assign cos[436]  =  16'b1100_0110_1101_0101;     //436pi/512
  assign sin[437]  =  16'b1110_0011_1001_0100;     //437pi/512
  assign cos[437]  =  16'b1100_0110_1010_1000;     //437pi/512
  assign sin[438]  =  16'b1110_0011_1110_1110;     //438pi/512
  assign cos[438]  =  16'b1100_0110_0111_1100;     //438pi/512
  assign sin[439]  =  16'b1110_0100_0100_1000;     //439pi/512
  assign cos[439]  =  16'b1100_0110_0101_0000;     //439pi/512
  assign sin[440]  =  16'b1110_0100_1010_0011;     //440pi/512
  assign cos[440]  =  16'b1100_0110_0010_0101;     //440pi/512
  assign sin[441]  =  16'b1110_0100_1111_1110;     //441pi/512
  assign cos[441]  =  16'b1100_0101_1111_1010;     //441pi/512
  assign sin[442]  =  16'b1110_0101_0101_1001;     //442pi/512
  assign cos[442]  =  16'b1100_0101_1101_0000;     //442pi/512
  assign sin[443]  =  16'b1110_0101_1011_0101;     //443pi/512
  assign cos[443]  =  16'b1100_0101_1010_0111;     //443pi/512
  assign sin[444]  =  16'b1110_0110_0001_0001;     //444pi/512
  assign cos[444]  =  16'b1100_0101_0111_1110;     //444pi/512
  assign sin[445]  =  16'b1110_0110_0110_1101;     //445pi/512
  assign cos[445]  =  16'b1100_0101_0101_0101;     //445pi/512
  assign sin[446]  =  16'b1110_0110_1100_1001;     //446pi/512
  assign cos[446]  =  16'b1100_0101_0010_1101;     //446pi/512
  assign sin[447]  =  16'b1110_0111_0010_0101;     //447pi/512
  assign cos[447]  =  16'b1100_0101_0000_0110;     //447pi/512
  assign sin[448]  =  16'b1110_0111_1000_0010;     //448pi/512
  assign cos[448]  =  16'b1100_0100_1101_1111;     //448pi/512
  assign sin[449]  =  16'b1110_0111_1101_1111;     //449pi/512
  assign cos[449]  =  16'b1100_0100_1011_1001;     //449pi/512
  assign sin[450]  =  16'b1110_1000_0011_1100;     //450pi/512
  assign cos[450]  =  16'b1100_0100_1001_0011;     //450pi/512
  assign sin[451]  =  16'b1110_1000_1001_1010;     //451pi/512
  assign cos[451]  =  16'b1100_0100_0110_1110;     //451pi/512
  assign sin[452]  =  16'b1110_1000_1111_0111;     //452pi/512
  assign cos[452]  =  16'b1100_0100_0100_1010;     //452pi/512
  assign sin[453]  =  16'b1110_1001_0101_0101;     //453pi/512
  assign cos[453]  =  16'b1100_0100_0010_0110;     //453pi/512
  assign sin[454]  =  16'b1110_1001_1011_0100;     //454pi/512
  assign cos[454]  =  16'b1100_0100_0000_0011;     //454pi/512
  assign sin[455]  =  16'b1110_1010_0001_0010;     //455pi/512
  assign cos[455]  =  16'b1100_0011_1110_0000;     //455pi/512
  assign sin[456]  =  16'b1110_1010_0111_0000;     //456pi/512
  assign cos[456]  =  16'b1100_0011_1011_1110;     //456pi/512
  assign sin[457]  =  16'b1110_1010_1100_1111;     //457pi/512
  assign cos[457]  =  16'b1100_0011_1001_1100;     //457pi/512
  assign sin[458]  =  16'b1110_1011_0010_1110;     //458pi/512
  assign cos[458]  =  16'b1100_0011_0111_1011;     //458pi/512
  assign sin[459]  =  16'b1110_1011_1000_1101;     //459pi/512
  assign cos[459]  =  16'b1100_0011_0101_1011;     //459pi/512
  assign sin[460]  =  16'b1110_1011_1110_1101;     //460pi/512
  assign cos[460]  =  16'b1100_0011_0011_1011;     //460pi/512
  assign sin[461]  =  16'b1110_1100_0100_1100;     //461pi/512
  assign cos[461]  =  16'b1100_0011_0001_1100;     //461pi/512
  assign sin[462]  =  16'b1110_1100_1010_1100;     //462pi/512
  assign cos[462]  =  16'b1100_0010_1111_1101;     //462pi/512
  assign sin[463]  =  16'b1110_1101_0000_1100;     //463pi/512
  assign cos[463]  =  16'b1100_0010_1101_1111;     //463pi/512
  assign sin[464]  =  16'b1110_1101_0110_1100;     //464pi/512
  assign cos[464]  =  16'b1100_0010_1100_0001;     //464pi/512
  assign sin[465]  =  16'b1110_1101_1100_1100;     //465pi/512
  assign cos[465]  =  16'b1100_0010_1010_0101;     //465pi/512
  assign sin[466]  =  16'b1110_1110_0010_1101;     //466pi/512
  assign cos[466]  =  16'b1100_0010_1000_1000;     //466pi/512
  assign sin[467]  =  16'b1110_1110_1000_1101;     //467pi/512
  assign cos[467]  =  16'b1100_0010_0110_1101;     //467pi/512
  assign sin[468]  =  16'b1110_1110_1110_1110;     //468pi/512
  assign cos[468]  =  16'b1100_0010_0101_0001;     //468pi/512
  assign sin[469]  =  16'b1110_1111_0100_1111;     //469pi/512
  assign cos[469]  =  16'b1100_0010_0011_0111;     //469pi/512
  assign sin[470]  =  16'b1110_1111_1011_0000;     //470pi/512
  assign cos[470]  =  16'b1100_0010_0001_1101;     //470pi/512
  assign sin[471]  =  16'b1111_0000_0001_0010;     //471pi/512
  assign cos[471]  =  16'b1100_0010_0000_0100;     //471pi/512
  assign sin[472]  =  16'b1111_0000_0111_0011;     //472pi/512
  assign cos[472]  =  16'b1100_0001_1110_1011;     //472pi/512
  assign sin[473]  =  16'b1111_0000_1101_0101;     //473pi/512
  assign cos[473]  =  16'b1100_0001_1101_0011;     //473pi/512
  assign sin[474]  =  16'b1111_0001_0011_0110;     //474pi/512
  assign cos[474]  =  16'b1100_0001_1011_1011;     //474pi/512
  assign sin[475]  =  16'b1111_0001_1001_1000;     //475pi/512
  assign cos[475]  =  16'b1100_0001_1010_0100;     //475pi/512
  assign sin[476]  =  16'b1111_0001_1111_1010;     //476pi/512
  assign cos[476]  =  16'b1100_0001_1000_1110;     //476pi/512
  assign sin[477]  =  16'b1111_0010_0101_1100;     //477pi/512
  assign cos[477]  =  16'b1100_0001_0111_1000;     //477pi/512
  assign sin[478]  =  16'b1111_0010_1011_1111;     //478pi/512
  assign cos[478]  =  16'b1100_0001_0110_0011;     //478pi/512
  assign sin[479]  =  16'b1111_0011_0010_0001;     //479pi/512
  assign cos[479]  =  16'b1100_0001_0100_1111;     //479pi/512
  assign sin[480]  =  16'b1111_0011_1000_0100;     //480pi/512
  assign cos[480]  =  16'b1100_0001_0011_1011;     //480pi/512
  assign sin[481]  =  16'b1111_0011_1110_0110;     //481pi/512
  assign cos[481]  =  16'b1100_0001_0010_1000;     //481pi/512
  assign sin[482]  =  16'b1111_0100_0100_1001;     //482pi/512
  assign cos[482]  =  16'b1100_0001_0001_0101;     //482pi/512
  assign sin[483]  =  16'b1111_0100_1010_1100;     //483pi/512
  assign cos[483]  =  16'b1100_0001_0000_0011;     //483pi/512
  assign sin[484]  =  16'b1111_0101_0000_1111;     //484pi/512
  assign cos[484]  =  16'b1100_0000_1111_0001;     //484pi/512
  assign sin[485]  =  16'b1111_0101_0111_0010;     //485pi/512
  assign cos[485]  =  16'b1100_0000_1110_0000;     //485pi/512
  assign sin[486]  =  16'b1111_0101_1101_0101;     //486pi/512
  assign cos[486]  =  16'b1100_0000_1101_0000;     //486pi/512
  assign sin[487]  =  16'b1111_0110_0011_1001;     //487pi/512
  assign cos[487]  =  16'b1100_0000_1100_0000;     //487pi/512
  assign sin[488]  =  16'b1111_0110_1001_1100;     //488pi/512
  assign cos[488]  =  16'b1100_0000_1011_0001;     //488pi/512
  assign sin[489]  =  16'b1111_0110_1111_1111;     //489pi/512
  assign cos[489]  =  16'b1100_0000_1010_0011;     //489pi/512
  assign sin[490]  =  16'b1111_0111_0110_0011;     //490pi/512
  assign cos[490]  =  16'b1100_0000_1001_0101;     //490pi/512
  assign sin[491]  =  16'b1111_0111_1100_0111;     //491pi/512
  assign cos[491]  =  16'b1100_0000_1000_1000;     //491pi/512
  assign sin[492]  =  16'b1111_1000_0010_1010;     //492pi/512
  assign cos[492]  =  16'b1100_0000_0111_1011;     //492pi/512
  assign sin[493]  =  16'b1111_1000_1000_1110;     //493pi/512
  assign cos[493]  =  16'b1100_0000_0110_1111;     //493pi/512
  assign sin[494]  =  16'b1111_1000_1111_0010;     //494pi/512
  assign cos[494]  =  16'b1100_0000_0110_0100;     //494pi/512
  assign sin[495]  =  16'b1111_1001_0101_0110;     //495pi/512
  assign cos[495]  =  16'b1100_0000_0101_1001;     //495pi/512
  assign sin[496]  =  16'b1111_1001_1011_1010;     //496pi/512
  assign cos[496]  =  16'b1100_0000_0100_1111;     //496pi/512
  assign sin[497]  =  16'b1111_1010_0001_1110;     //497pi/512
  assign cos[497]  =  16'b1100_0000_0100_0101;     //497pi/512
  assign sin[498]  =  16'b1111_1010_1000_0010;     //498pi/512
  assign cos[498]  =  16'b1100_0000_0011_1100;     //498pi/512
  assign sin[499]  =  16'b1111_1010_1110_0110;     //499pi/512
  assign cos[499]  =  16'b1100_0000_0011_0100;     //499pi/512
  assign sin[500]  =  16'b1111_1011_0100_1011;     //500pi/512
  assign cos[500]  =  16'b1100_0000_0010_1100;     //500pi/512
  assign sin[501]  =  16'b1111_1011_1010_1111;     //501pi/512
  assign cos[501]  =  16'b1100_0000_0010_0101;     //501pi/512
  assign sin[502]  =  16'b1111_1100_0001_0011;     //502pi/512
  assign cos[502]  =  16'b1100_0000_0001_1111;     //502pi/512
  assign sin[503]  =  16'b1111_1100_0111_1000;     //503pi/512
  assign cos[503]  =  16'b1100_0000_0001_1001;     //503pi/512
  assign sin[504]  =  16'b1111_1100_1101_1100;     //504pi/512
  assign cos[504]  =  16'b1100_0000_0001_0100;     //504pi/512
  assign sin[505]  =  16'b1111_1101_0100_0000;     //505pi/512
  assign cos[505]  =  16'b1100_0000_0000_1111;     //505pi/512
  assign sin[506]  =  16'b1111_1101_1010_0101;     //506pi/512
  assign cos[506]  =  16'b1100_0000_0000_1011;     //506pi/512
  assign sin[507]  =  16'b1111_1110_0000_1001;     //507pi/512
  assign cos[507]  =  16'b1100_0000_0000_1000;     //507pi/512
  assign sin[508]  =  16'b1111_1110_0110_1110;     //508pi/512
  assign cos[508]  =  16'b1100_0000_0000_0101;     //508pi/512
  assign sin[509]  =  16'b1111_1110_1101_0010;     //509pi/512
  assign cos[509]  =  16'b1100_0000_0000_0011;     //509pi/512
  assign sin[510]  =  16'b1111_1111_0011_0111;     //510pi/512
  assign cos[510]  =  16'b1100_0000_0000_0001;     //510pi/512
  assign sin[511]  =  16'b1111_1111_1001_1011;     //511pi/512
  assign cos[511]  =  16'b1100_0000_0000_0000;     //511pi/512

endmodule