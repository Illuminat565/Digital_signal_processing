module  tw_factor_for_6th #(parameter stage_FFT = 2, SIZE =10, word_length_tw = 14) (
    input            clk,
    input            en_rd, 
    input   [stage_FFT-2:0]   rd_ptr_angle,

    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );


reg signed [word_length_tw-1:0]  cos  [31:0];
reg signed [word_length_tw-1:0]  sin  [31:0];


//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd  ) begin
                  cos_data           <= cos   [rd_ptr_angle];
                  sin_data           <= sin   [rd_ptr_angle];
             end 
        end

//--------------------------------handle read tw factor------------------------------

initial begin
   sin[0]  =  14'b00000000000000;     //0pi/256
   cos[0]  =  14'b01000000000000;     //0pi/256
   sin[1]  =  14'b11111001101111;     //8pi/256
   cos[1]  =  14'b00111111101100;     //8pi/256
   sin[2]  =  14'b11110011100001;     //16pi/256
   cos[2]  =  14'b00111110110001;     //16pi/256
   sin[3]  =  14'b11101101011011;     //24pi/256
   cos[3]  =  14'b00111101001111;     //24pi/256
   sin[4]  =  14'b11100111100001;     //32pi/256
   cos[4]  =  14'b00111011001000;     //32pi/256
   sin[5]  =  14'b11100001110101;     //40pi/256
   cos[5]  =  14'b00111000011100;     //40pi/256
   sin[6]  =  14'b11011100011100;     //48pi/256
   cos[6]  =  14'b00110101001101;     //48pi/256
   sin[7]  =  14'b11010111011010;     //56pi/256
   cos[7]  =  14'b00110001011110;     //56pi/256
   sin[8]  =  14'b11010010110000;     //64pi/256
   cos[8]  =  14'b00101101010000;     //64pi/256
   sin[9]  =  14'b11001110100010;     //72pi/256
   cos[9]  =  14'b00101000100110;     //72pi/256
   sin[10]  =  14'b11001010110010;     //80pi/256
   cos[10]  =  14'b00100011100011;     //80pi/256
   sin[11]  =  14'b11000111100100;     //88pi/256
   cos[11]  =  14'b00011110001010;     //88pi/256
   sin[12]  =  14'b11000100111000;     //96pi/256
   cos[12]  =  14'b00011000011111;     //96pi/256
   sin[13]  =  14'b11000010110000;     //104pi/256
   cos[13]  =  14'b00010010100101;     //104pi/256
   sin[14]  =  14'b11000001001111;     //112pi/256
   cos[14]  =  14'b00001100011111;     //112pi/256
   sin[15]  =  14'b11000000010100;     //120pi/256
   cos[15]  =  14'b00000110010001;     //120pi/256
   sin[16]  =  14'b11000000000000;     //128pi/256
   cos[16]  =  14'b00000000000000;     //128pi/256
   sin[17]  =  14'b11000000010100;     //136pi/256
   cos[17]  =  14'b11111001101111;     //136pi/256
   sin[18]  =  14'b11000001001111;     //144pi/256
   cos[18]  =  14'b11110011100001;     //144pi/256
   sin[19]  =  14'b11000010110000;     //152pi/256
   cos[19]  =  14'b11101101011011;     //152pi/256
   sin[20]  =  14'b11000100111000;     //160pi/256
   cos[20]  =  14'b11100111100001;     //160pi/256
   sin[21]  =  14'b11000111100100;     //168pi/256
   cos[21]  =  14'b11100001110101;     //168pi/256
   sin[22]  =  14'b11001010110010;     //176pi/256
   cos[22]  =  14'b11011100011100;     //176pi/256
   sin[23]  =  14'b11001110100010;     //184pi/256
   cos[23]  =  14'b11010111011010;     //184pi/256
   sin[24]  =  14'b11010010110000;     //192pi/256
   cos[24]  =  14'b11010010110000;     //192pi/256
   sin[25]  =  14'b11010111011010;     //200pi/256
   cos[25]  =  14'b11001110100010;     //200pi/256
   sin[26]  =  14'b11011100011100;     //208pi/256
   cos[26]  =  14'b11001010110010;     //208pi/256
   sin[27]  =  14'b11100001110101;     //216pi/256
   cos[27]  =  14'b11000111100100;     //216pi/256
   sin[28]  =  14'b11100111100001;     //224pi/256
   cos[28]  =  14'b11000100111000;     //224pi/256
   sin[29]  =  14'b11101101011011;     //232pi/256
   cos[29]  =  14'b11000010110000;     //232pi/256
   sin[30]  =  14'b11110011100001;     //240pi/256
   cos[30]  =  14'b11000001001111;     //240pi/256
   sin[31]  =  14'b11111001101111;     //248pi/256
   cos[31]  =  14'b11000000010100;     //248pi/256
end
endmodule