module  M_TWIDLE_13_B_0_10_v  #(parameter SIZE = 10, word_length_tw = 13) (
    input            clk,
    input            en_rd,
    input   [10:0]   rd_ptr_angle,
    input            en_modf,
    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );
reg signed [word_length_tw-1:0]  cos    [511:0];
reg signed [word_length_tw-1:0]  sin    [511:0];
reg signed [word_length_tw-1:0]  m_cos  [511:0];
reg signed [word_length_tw-1:0]  m_sin  [511:0];
reg signed [word_length_tw-1:0]  cos_temp;
reg signed [word_length_tw-1:0]  sin_temp;
reg signed [word_length_tw-1:0]  m_cos_temp;
reg signed [word_length_tw-1:0]  m_sin_temp;
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & ~ en_modf) begin
                  cos_temp           <= cos   [rd_ptr_angle];
                  sin_temp           <= sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & en_modf) begin
                  m_cos_temp           <= m_cos   [rd_ptr_angle];
                  m_sin_temp           <= m_sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(*) begin 
             if (en_modf) begin
                  cos_data           <= m_cos_temp;
                  sin_data           <= m_sin_temp;
             end else begin
                  cos_data           <= cos_temp;
                  sin_data           <= sin_temp;
             end 
        end
initial begin
   sin[0]  =  13'b0000000000000;     //0pi/512
   cos[0]  =  13'b0100000000000;     //0pi/512
   sin[1]  =  13'b1111111110011;     //1pi/512
   cos[1]  =  13'b0011111111111;     //1pi/512
   sin[2]  =  13'b1111111100111;     //2pi/512
   cos[2]  =  13'b0011111111111;     //2pi/512
   sin[3]  =  13'b1111111011010;     //3pi/512
   cos[3]  =  13'b0011111111111;     //3pi/512
   sin[4]  =  13'b1111111001110;     //4pi/512
   cos[4]  =  13'b0011111111111;     //4pi/512
   sin[5]  =  13'b1111111000001;     //5pi/512
   cos[5]  =  13'b0011111111111;     //5pi/512
   sin[6]  =  13'b1111110110101;     //6pi/512
   cos[6]  =  13'b0011111111110;     //6pi/512
   sin[7]  =  13'b1111110101000;     //7pi/512
   cos[7]  =  13'b0011111111110;     //7pi/512
   sin[8]  =  13'b1111110011100;     //8pi/512
   cos[8]  =  13'b0011111111101;     //8pi/512
   sin[9]  =  13'b1111110001111;     //9pi/512
   cos[9]  =  13'b0011111111100;     //9pi/512
   sin[10]  =  13'b1111110000010;     //10pi/512
   cos[10]  =  13'b0011111111100;     //10pi/512
   sin[11]  =  13'b1111101110110;     //11pi/512
   cos[11]  =  13'b0011111111011;     //11pi/512
   sin[12]  =  13'b1111101101001;     //12pi/512
   cos[12]  =  13'b0011111111010;     //12pi/512
   sin[13]  =  13'b1111101011101;     //13pi/512
   cos[13]  =  13'b0011111111001;     //13pi/512
   sin[14]  =  13'b1111101010000;     //14pi/512
   cos[14]  =  13'b0011111111000;     //14pi/512
   sin[15]  =  13'b1111101000100;     //15pi/512
   cos[15]  =  13'b0011111110111;     //15pi/512
   sin[16]  =  13'b1111100110111;     //16pi/512
   cos[16]  =  13'b0011111110110;     //16pi/512
   sin[17]  =  13'b1111100101011;     //17pi/512
   cos[17]  =  13'b0011111110100;     //17pi/512
   sin[18]  =  13'b1111100011110;     //18pi/512
   cos[18]  =  13'b0011111110011;     //18pi/512
   sin[19]  =  13'b1111100010010;     //19pi/512
   cos[19]  =  13'b0011111110010;     //19pi/512
   sin[20]  =  13'b1111100000101;     //20pi/512
   cos[20]  =  13'b0011111110000;     //20pi/512
   sin[21]  =  13'b1111011111001;     //21pi/512
   cos[21]  =  13'b0011111101111;     //21pi/512
   sin[22]  =  13'b1111011101100;     //22pi/512
   cos[22]  =  13'b0011111101101;     //22pi/512
   sin[23]  =  13'b1111011100000;     //23pi/512
   cos[23]  =  13'b0011111101011;     //23pi/512
   sin[24]  =  13'b1111011010011;     //24pi/512
   cos[24]  =  13'b0011111101001;     //24pi/512
   sin[25]  =  13'b1111011000111;     //25pi/512
   cos[25]  =  13'b0011111100111;     //25pi/512
   sin[26]  =  13'b1111010111011;     //26pi/512
   cos[26]  =  13'b0011111100101;     //26pi/512
   sin[27]  =  13'b1111010101110;     //27pi/512
   cos[27]  =  13'b0011111100011;     //27pi/512
   sin[28]  =  13'b1111010100010;     //28pi/512
   cos[28]  =  13'b0011111100001;     //28pi/512
   sin[29]  =  13'b1111010010101;     //29pi/512
   cos[29]  =  13'b0011111011111;     //29pi/512
   sin[30]  =  13'b1111010001001;     //30pi/512
   cos[30]  =  13'b0011111011101;     //30pi/512
   sin[31]  =  13'b1111001111101;     //31pi/512
   cos[31]  =  13'b0011111011011;     //31pi/512
   sin[32]  =  13'b1111001110000;     //32pi/512
   cos[32]  =  13'b0011111011000;     //32pi/512
   sin[33]  =  13'b1111001100100;     //33pi/512
   cos[33]  =  13'b0011111010110;     //33pi/512
   sin[34]  =  13'b1111001011000;     //34pi/512
   cos[34]  =  13'b0011111010011;     //34pi/512
   sin[35]  =  13'b1111001001100;     //35pi/512
   cos[35]  =  13'b0011111010000;     //35pi/512
   sin[36]  =  13'b1111000111111;     //36pi/512
   cos[36]  =  13'b0011111001110;     //36pi/512
   sin[37]  =  13'b1111000110011;     //37pi/512
   cos[37]  =  13'b0011111001011;     //37pi/512
   sin[38]  =  13'b1111000100111;     //38pi/512
   cos[38]  =  13'b0011111001000;     //38pi/512
   sin[39]  =  13'b1111000011011;     //39pi/512
   cos[39]  =  13'b0011111000101;     //39pi/512
   sin[40]  =  13'b1111000001110;     //40pi/512
   cos[40]  =  13'b0011111000010;     //40pi/512
   sin[41]  =  13'b1111000000010;     //41pi/512
   cos[41]  =  13'b0011110111111;     //41pi/512
   sin[42]  =  13'b1110111110110;     //42pi/512
   cos[42]  =  13'b0011110111100;     //42pi/512
   sin[43]  =  13'b1110111101010;     //43pi/512
   cos[43]  =  13'b0011110111001;     //43pi/512
   sin[44]  =  13'b1110111011110;     //44pi/512
   cos[44]  =  13'b0011110110101;     //44pi/512
   sin[45]  =  13'b1110111010010;     //45pi/512
   cos[45]  =  13'b0011110110010;     //45pi/512
   sin[46]  =  13'b1110111000110;     //46pi/512
   cos[46]  =  13'b0011110101110;     //46pi/512
   sin[47]  =  13'b1110110111010;     //47pi/512
   cos[47]  =  13'b0011110101011;     //47pi/512
   sin[48]  =  13'b1110110101101;     //48pi/512
   cos[48]  =  13'b0011110100111;     //48pi/512
   sin[49]  =  13'b1110110100001;     //49pi/512
   cos[49]  =  13'b0011110100100;     //49pi/512
   sin[50]  =  13'b1110110010101;     //50pi/512
   cos[50]  =  13'b0011110100000;     //50pi/512
   sin[51]  =  13'b1110110001010;     //51pi/512
   cos[51]  =  13'b0011110011100;     //51pi/512
   sin[52]  =  13'b1110101111110;     //52pi/512
   cos[52]  =  13'b0011110011000;     //52pi/512
   sin[53]  =  13'b1110101110010;     //53pi/512
   cos[53]  =  13'b0011110010100;     //53pi/512
   sin[54]  =  13'b1110101100110;     //54pi/512
   cos[54]  =  13'b0011110010000;     //54pi/512
   sin[55]  =  13'b1110101011010;     //55pi/512
   cos[55]  =  13'b0011110001100;     //55pi/512
   sin[56]  =  13'b1110101001110;     //56pi/512
   cos[56]  =  13'b0011110001000;     //56pi/512
   sin[57]  =  13'b1110101000010;     //57pi/512
   cos[57]  =  13'b0011110000100;     //57pi/512
   sin[58]  =  13'b1110100110110;     //58pi/512
   cos[58]  =  13'b0011101111111;     //58pi/512
   sin[59]  =  13'b1110100101011;     //59pi/512
   cos[59]  =  13'b0011101111011;     //59pi/512
   sin[60]  =  13'b1110100011111;     //60pi/512
   cos[60]  =  13'b0011101110110;     //60pi/512
   sin[61]  =  13'b1110100010011;     //61pi/512
   cos[61]  =  13'b0011101110010;     //61pi/512
   sin[62]  =  13'b1110100001000;     //62pi/512
   cos[62]  =  13'b0011101101101;     //62pi/512
   sin[63]  =  13'b1110011111100;     //63pi/512
   cos[63]  =  13'b0011101101000;     //63pi/512
   sin[64]  =  13'b1110011110000;     //64pi/512
   cos[64]  =  13'b0011101100100;     //64pi/512
   sin[65]  =  13'b1110011100101;     //65pi/512
   cos[65]  =  13'b0011101011111;     //65pi/512
   sin[66]  =  13'b1110011011001;     //66pi/512
   cos[66]  =  13'b0011101011010;     //66pi/512
   sin[67]  =  13'b1110011001110;     //67pi/512
   cos[67]  =  13'b0011101010101;     //67pi/512
   sin[68]  =  13'b1110011000010;     //68pi/512
   cos[68]  =  13'b0011101010000;     //68pi/512
   sin[69]  =  13'b1110010110111;     //69pi/512
   cos[69]  =  13'b0011101001011;     //69pi/512
   sin[70]  =  13'b1110010101011;     //70pi/512
   cos[70]  =  13'b0011101000101;     //70pi/512
   sin[71]  =  13'b1110010100000;     //71pi/512
   cos[71]  =  13'b0011101000000;     //71pi/512
   sin[72]  =  13'b1110010010100;     //72pi/512
   cos[72]  =  13'b0011100111011;     //72pi/512
   sin[73]  =  13'b1110010001001;     //73pi/512
   cos[73]  =  13'b0011100110101;     //73pi/512
   sin[74]  =  13'b1110001111110;     //74pi/512
   cos[74]  =  13'b0011100110000;     //74pi/512
   sin[75]  =  13'b1110001110010;     //75pi/512
   cos[75]  =  13'b0011100101010;     //75pi/512
   sin[76]  =  13'b1110001100111;     //76pi/512
   cos[76]  =  13'b0011100100101;     //76pi/512
   sin[77]  =  13'b1110001011100;     //77pi/512
   cos[77]  =  13'b0011100011111;     //77pi/512
   sin[78]  =  13'b1110001010001;     //78pi/512
   cos[78]  =  13'b0011100011001;     //78pi/512
   sin[79]  =  13'b1110001000110;     //79pi/512
   cos[79]  =  13'b0011100010100;     //79pi/512
   sin[80]  =  13'b1110000111011;     //80pi/512
   cos[80]  =  13'b0011100001110;     //80pi/512
   sin[81]  =  13'b1110000110000;     //81pi/512
   cos[81]  =  13'b0011100001000;     //81pi/512
   sin[82]  =  13'b1110000100100;     //82pi/512
   cos[82]  =  13'b0011100000010;     //82pi/512
   sin[83]  =  13'b1110000011001;     //83pi/512
   cos[83]  =  13'b0011011111100;     //83pi/512
   sin[84]  =  13'b1110000001111;     //84pi/512
   cos[84]  =  13'b0011011110101;     //84pi/512
   sin[85]  =  13'b1110000000100;     //85pi/512
   cos[85]  =  13'b0011011101111;     //85pi/512
   sin[86]  =  13'b1101111111001;     //86pi/512
   cos[86]  =  13'b0011011101001;     //86pi/512
   sin[87]  =  13'b1101111101110;     //87pi/512
   cos[87]  =  13'b0011011100011;     //87pi/512
   sin[88]  =  13'b1101111100011;     //88pi/512
   cos[88]  =  13'b0011011011100;     //88pi/512
   sin[89]  =  13'b1101111011000;     //89pi/512
   cos[89]  =  13'b0011011010110;     //89pi/512
   sin[90]  =  13'b1101111001110;     //90pi/512
   cos[90]  =  13'b0011011001111;     //90pi/512
   sin[91]  =  13'b1101111000011;     //91pi/512
   cos[91]  =  13'b0011011001000;     //91pi/512
   sin[92]  =  13'b1101110111000;     //92pi/512
   cos[92]  =  13'b0011011000010;     //92pi/512
   sin[93]  =  13'b1101110101110;     //93pi/512
   cos[93]  =  13'b0011010111011;     //93pi/512
   sin[94]  =  13'b1101110100011;     //94pi/512
   cos[94]  =  13'b0011010110100;     //94pi/512
   sin[95]  =  13'b1101110011001;     //95pi/512
   cos[95]  =  13'b0011010101101;     //95pi/512
   sin[96]  =  13'b1101110001110;     //96pi/512
   cos[96]  =  13'b0011010100110;     //96pi/512
   sin[97]  =  13'b1101110000100;     //97pi/512
   cos[97]  =  13'b0011010011111;     //97pi/512
   sin[98]  =  13'b1101101111001;     //98pi/512
   cos[98]  =  13'b0011010011000;     //98pi/512
   sin[99]  =  13'b1101101101111;     //99pi/512
   cos[99]  =  13'b0011010010001;     //99pi/512
   sin[100]  =  13'b1101101100101;     //100pi/512
   cos[100]  =  13'b0011010001010;     //100pi/512
   sin[101]  =  13'b1101101011010;     //101pi/512
   cos[101]  =  13'b0011010000011;     //101pi/512
   sin[102]  =  13'b1101101010000;     //102pi/512
   cos[102]  =  13'b0011001111011;     //102pi/512
   sin[103]  =  13'b1101101000110;     //103pi/512
   cos[103]  =  13'b0011001110100;     //103pi/512
   sin[104]  =  13'b1101100111100;     //104pi/512
   cos[104]  =  13'b0011001101100;     //104pi/512
   sin[105]  =  13'b1101100110010;     //105pi/512
   cos[105]  =  13'b0011001100101;     //105pi/512
   sin[106]  =  13'b1101100101000;     //106pi/512
   cos[106]  =  13'b0011001011101;     //106pi/512
   sin[107]  =  13'b1101100011110;     //107pi/512
   cos[107]  =  13'b0011001010110;     //107pi/512
   sin[108]  =  13'b1101100010100;     //108pi/512
   cos[108]  =  13'b0011001001110;     //108pi/512
   sin[109]  =  13'b1101100001010;     //109pi/512
   cos[109]  =  13'b0011001000110;     //109pi/512
   sin[110]  =  13'b1101100000000;     //110pi/512
   cos[110]  =  13'b0011000111110;     //110pi/512
   sin[111]  =  13'b1101011110111;     //111pi/512
   cos[111]  =  13'b0011000110111;     //111pi/512
   sin[112]  =  13'b1101011101101;     //112pi/512
   cos[112]  =  13'b0011000101111;     //112pi/512
   sin[113]  =  13'b1101011100011;     //113pi/512
   cos[113]  =  13'b0011000100111;     //113pi/512
   sin[114]  =  13'b1101011011001;     //114pi/512
   cos[114]  =  13'b0011000011111;     //114pi/512
   sin[115]  =  13'b1101011010000;     //115pi/512
   cos[115]  =  13'b0011000010110;     //115pi/512
   sin[116]  =  13'b1101011000110;     //116pi/512
   cos[116]  =  13'b0011000001110;     //116pi/512
   sin[117]  =  13'b1101010111101;     //117pi/512
   cos[117]  =  13'b0011000000110;     //117pi/512
   sin[118]  =  13'b1101010110011;     //118pi/512
   cos[118]  =  13'b0010111111110;     //118pi/512
   sin[119]  =  13'b1101010101010;     //119pi/512
   cos[119]  =  13'b0010111110101;     //119pi/512
   sin[120]  =  13'b1101010100001;     //120pi/512
   cos[120]  =  13'b0010111101101;     //120pi/512
   sin[121]  =  13'b1101010010111;     //121pi/512
   cos[121]  =  13'b0010111100101;     //121pi/512
   sin[122]  =  13'b1101010001110;     //122pi/512
   cos[122]  =  13'b0010111011100;     //122pi/512
   sin[123]  =  13'b1101010000101;     //123pi/512
   cos[123]  =  13'b0010111010011;     //123pi/512
   sin[124]  =  13'b1101001111100;     //124pi/512
   cos[124]  =  13'b0010111001011;     //124pi/512
   sin[125]  =  13'b1101001110011;     //125pi/512
   cos[125]  =  13'b0010111000010;     //125pi/512
   sin[126]  =  13'b1101001101010;     //126pi/512
   cos[126]  =  13'b0010110111001;     //126pi/512
   sin[127]  =  13'b1101001100001;     //127pi/512
   cos[127]  =  13'b0010110110001;     //127pi/512
   sin[128]  =  13'b1101001011000;     //128pi/512
   cos[128]  =  13'b0010110101000;     //128pi/512
   sin[129]  =  13'b1101001001111;     //129pi/512
   cos[129]  =  13'b0010110011111;     //129pi/512
   sin[130]  =  13'b1101001000110;     //130pi/512
   cos[130]  =  13'b0010110010110;     //130pi/512
   sin[131]  =  13'b1101000111101;     //131pi/512
   cos[131]  =  13'b0010110001101;     //131pi/512
   sin[132]  =  13'b1101000110101;     //132pi/512
   cos[132]  =  13'b0010110000100;     //132pi/512
   sin[133]  =  13'b1101000101100;     //133pi/512
   cos[133]  =  13'b0010101111011;     //133pi/512
   sin[134]  =  13'b1101000100100;     //134pi/512
   cos[134]  =  13'b0010101110001;     //134pi/512
   sin[135]  =  13'b1101000011011;     //135pi/512
   cos[135]  =  13'b0010101101000;     //135pi/512
   sin[136]  =  13'b1101000010011;     //136pi/512
   cos[136]  =  13'b0010101011111;     //136pi/512
   sin[137]  =  13'b1101000001010;     //137pi/512
   cos[137]  =  13'b0010101010110;     //137pi/512
   sin[138]  =  13'b1101000000010;     //138pi/512
   cos[138]  =  13'b0010101001100;     //138pi/512
   sin[139]  =  13'b1100111111001;     //139pi/512
   cos[139]  =  13'b0010101000011;     //139pi/512
   sin[140]  =  13'b1100111110001;     //140pi/512
   cos[140]  =  13'b0010100111001;     //140pi/512
   sin[141]  =  13'b1100111101001;     //141pi/512
   cos[141]  =  13'b0010100110000;     //141pi/512
   sin[142]  =  13'b1100111100001;     //142pi/512
   cos[142]  =  13'b0010100100110;     //142pi/512
   sin[143]  =  13'b1100111011001;     //143pi/512
   cos[143]  =  13'b0010100011100;     //143pi/512
   sin[144]  =  13'b1100111010001;     //144pi/512
   cos[144]  =  13'b0010100010011;     //144pi/512
   sin[145]  =  13'b1100111001001;     //145pi/512
   cos[145]  =  13'b0010100001001;     //145pi/512
   sin[146]  =  13'b1100111000001;     //146pi/512
   cos[146]  =  13'b0010011111111;     //146pi/512
   sin[147]  =  13'b1100110111001;     //147pi/512
   cos[147]  =  13'b0010011110101;     //147pi/512
   sin[148]  =  13'b1100110110001;     //148pi/512
   cos[148]  =  13'b0010011101011;     //148pi/512
   sin[149]  =  13'b1100110101010;     //149pi/512
   cos[149]  =  13'b0010011100010;     //149pi/512
   sin[150]  =  13'b1100110100010;     //150pi/512
   cos[150]  =  13'b0010011011000;     //150pi/512
   sin[151]  =  13'b1100110011011;     //151pi/512
   cos[151]  =  13'b0010011001110;     //151pi/512
   sin[152]  =  13'b1100110010011;     //152pi/512
   cos[152]  =  13'b0010011000011;     //152pi/512
   sin[153]  =  13'b1100110001100;     //153pi/512
   cos[153]  =  13'b0010010111001;     //153pi/512
   sin[154]  =  13'b1100110000100;     //154pi/512
   cos[154]  =  13'b0010010101111;     //154pi/512
   sin[155]  =  13'b1100101111101;     //155pi/512
   cos[155]  =  13'b0010010100101;     //155pi/512
   sin[156]  =  13'b1100101110110;     //156pi/512
   cos[156]  =  13'b0010010011011;     //156pi/512
   sin[157]  =  13'b1100101101110;     //157pi/512
   cos[157]  =  13'b0010010010000;     //157pi/512
   sin[158]  =  13'b1100101100111;     //158pi/512
   cos[158]  =  13'b0010010000110;     //158pi/512
   sin[159]  =  13'b1100101100000;     //159pi/512
   cos[159]  =  13'b0010001111100;     //159pi/512
   sin[160]  =  13'b1100101011001;     //160pi/512
   cos[160]  =  13'b0010001110001;     //160pi/512
   sin[161]  =  13'b1100101010010;     //161pi/512
   cos[161]  =  13'b0010001100111;     //161pi/512
   sin[162]  =  13'b1100101001011;     //162pi/512
   cos[162]  =  13'b0010001011100;     //162pi/512
   sin[163]  =  13'b1100101000100;     //163pi/512
   cos[163]  =  13'b0010001010010;     //163pi/512
   sin[164]  =  13'b1100100111110;     //164pi/512
   cos[164]  =  13'b0010001000111;     //164pi/512
   sin[165]  =  13'b1100100110111;     //165pi/512
   cos[165]  =  13'b0010000111101;     //165pi/512
   sin[166]  =  13'b1100100110000;     //166pi/512
   cos[166]  =  13'b0010000110010;     //166pi/512
   sin[167]  =  13'b1100100101010;     //167pi/512
   cos[167]  =  13'b0010000100111;     //167pi/512
   sin[168]  =  13'b1100100100011;     //168pi/512
   cos[168]  =  13'b0010000011100;     //168pi/512
   sin[169]  =  13'b1100100011101;     //169pi/512
   cos[169]  =  13'b0010000010010;     //169pi/512
   sin[170]  =  13'b1100100010111;     //170pi/512
   cos[170]  =  13'b0010000000111;     //170pi/512
   sin[171]  =  13'b1100100010000;     //171pi/512
   cos[171]  =  13'b0001111111100;     //171pi/512
   sin[172]  =  13'b1100100001010;     //172pi/512
   cos[172]  =  13'b0001111110001;     //172pi/512
   sin[173]  =  13'b1100100000100;     //173pi/512
   cos[173]  =  13'b0001111100110;     //173pi/512
   sin[174]  =  13'b1100011111110;     //174pi/512
   cos[174]  =  13'b0001111011011;     //174pi/512
   sin[175]  =  13'b1100011111000;     //175pi/512
   cos[175]  =  13'b0001111010000;     //175pi/512
   sin[176]  =  13'b1100011110010;     //176pi/512
   cos[176]  =  13'b0001111000101;     //176pi/512
   sin[177]  =  13'b1100011101100;     //177pi/512
   cos[177]  =  13'b0001110111010;     //177pi/512
   sin[178]  =  13'b1100011100110;     //178pi/512
   cos[178]  =  13'b0001110101111;     //178pi/512
   sin[179]  =  13'b1100011100000;     //179pi/512
   cos[179]  =  13'b0001110100100;     //179pi/512
   sin[180]  =  13'b1100011011011;     //180pi/512
   cos[180]  =  13'b0001110011000;     //180pi/512
   sin[181]  =  13'b1100011010101;     //181pi/512
   cos[181]  =  13'b0001110001101;     //181pi/512
   sin[182]  =  13'b1100011010000;     //182pi/512
   cos[182]  =  13'b0001110000010;     //182pi/512
   sin[183]  =  13'b1100011001010;     //183pi/512
   cos[183]  =  13'b0001101110110;     //183pi/512
   sin[184]  =  13'b1100011000101;     //184pi/512
   cos[184]  =  13'b0001101101011;     //184pi/512
   sin[185]  =  13'b1100010111111;     //185pi/512
   cos[185]  =  13'b0001101100000;     //185pi/512
   sin[186]  =  13'b1100010111010;     //186pi/512
   cos[186]  =  13'b0001101010100;     //186pi/512
   sin[187]  =  13'b1100010110101;     //187pi/512
   cos[187]  =  13'b0001101001001;     //187pi/512
   sin[188]  =  13'b1100010110000;     //188pi/512
   cos[188]  =  13'b0001100111101;     //188pi/512
   sin[189]  =  13'b1100010101011;     //189pi/512
   cos[189]  =  13'b0001100110010;     //189pi/512
   sin[190]  =  13'b1100010100110;     //190pi/512
   cos[190]  =  13'b0001100100110;     //190pi/512
   sin[191]  =  13'b1100010100001;     //191pi/512
   cos[191]  =  13'b0001100011011;     //191pi/512
   sin[192]  =  13'b1100010011100;     //192pi/512
   cos[192]  =  13'b0001100001111;     //192pi/512
   sin[193]  =  13'b1100010010111;     //193pi/512
   cos[193]  =  13'b0001100000100;     //193pi/512
   sin[194]  =  13'b1100010010010;     //194pi/512
   cos[194]  =  13'b0001011111000;     //194pi/512
   sin[195]  =  13'b1100010001110;     //195pi/512
   cos[195]  =  13'b0001011101100;     //195pi/512
   sin[196]  =  13'b1100010001001;     //196pi/512
   cos[196]  =  13'b0001011100001;     //196pi/512
   sin[197]  =  13'b1100010000101;     //197pi/512
   cos[197]  =  13'b0001011010101;     //197pi/512
   sin[198]  =  13'b1100010000000;     //198pi/512
   cos[198]  =  13'b0001011001001;     //198pi/512
   sin[199]  =  13'b1100001111100;     //199pi/512
   cos[199]  =  13'b0001010111101;     //199pi/512
   sin[200]  =  13'b1100001111000;     //200pi/512
   cos[200]  =  13'b0001010110001;     //200pi/512
   sin[201]  =  13'b1100001110100;     //201pi/512
   cos[201]  =  13'b0001010100110;     //201pi/512
   sin[202]  =  13'b1100001101111;     //202pi/512
   cos[202]  =  13'b0001010011010;     //202pi/512
   sin[203]  =  13'b1100001101011;     //203pi/512
   cos[203]  =  13'b0001010001110;     //203pi/512
   sin[204]  =  13'b1100001100111;     //204pi/512
   cos[204]  =  13'b0001010000010;     //204pi/512
   sin[205]  =  13'b1100001100011;     //205pi/512
   cos[205]  =  13'b0001001110110;     //205pi/512
   sin[206]  =  13'b1100001100000;     //206pi/512
   cos[206]  =  13'b0001001101010;     //206pi/512
   sin[207]  =  13'b1100001011100;     //207pi/512
   cos[207]  =  13'b0001001011110;     //207pi/512
   sin[208]  =  13'b1100001011000;     //208pi/512
   cos[208]  =  13'b0001001010010;     //208pi/512
   sin[209]  =  13'b1100001010101;     //209pi/512
   cos[209]  =  13'b0001001000110;     //209pi/512
   sin[210]  =  13'b1100001010001;     //210pi/512
   cos[210]  =  13'b0001000111010;     //210pi/512
   sin[211]  =  13'b1100001001110;     //211pi/512
   cos[211]  =  13'b0001000101110;     //211pi/512
   sin[212]  =  13'b1100001001010;     //212pi/512
   cos[212]  =  13'b0001000100010;     //212pi/512
   sin[213]  =  13'b1100001000111;     //213pi/512
   cos[213]  =  13'b0001000010110;     //213pi/512
   sin[214]  =  13'b1100001000100;     //214pi/512
   cos[214]  =  13'b0001000001001;     //214pi/512
   sin[215]  =  13'b1100001000000;     //215pi/512
   cos[215]  =  13'b0000111111101;     //215pi/512
   sin[216]  =  13'b1100000111101;     //216pi/512
   cos[216]  =  13'b0000111110001;     //216pi/512
   sin[217]  =  13'b1100000111010;     //217pi/512
   cos[217]  =  13'b0000111100101;     //217pi/512
   sin[218]  =  13'b1100000110111;     //218pi/512
   cos[218]  =  13'b0000111011001;     //218pi/512
   sin[219]  =  13'b1100000110101;     //219pi/512
   cos[219]  =  13'b0000111001100;     //219pi/512
   sin[220]  =  13'b1100000110010;     //220pi/512
   cos[220]  =  13'b0000111000000;     //220pi/512
   sin[221]  =  13'b1100000101111;     //221pi/512
   cos[221]  =  13'b0000110110100;     //221pi/512
   sin[222]  =  13'b1100000101100;     //222pi/512
   cos[222]  =  13'b0000110101000;     //222pi/512
   sin[223]  =  13'b1100000101010;     //223pi/512
   cos[223]  =  13'b0000110011011;     //223pi/512
   sin[224]  =  13'b1100000100111;     //224pi/512
   cos[224]  =  13'b0000110001111;     //224pi/512
   sin[225]  =  13'b1100000100101;     //225pi/512
   cos[225]  =  13'b0000110000011;     //225pi/512
   sin[226]  =  13'b1100000100011;     //226pi/512
   cos[226]  =  13'b0000101110110;     //226pi/512
   sin[227]  =  13'b1100000100000;     //227pi/512
   cos[227]  =  13'b0000101101010;     //227pi/512
   sin[228]  =  13'b1100000011110;     //228pi/512
   cos[228]  =  13'b0000101011110;     //228pi/512
   sin[229]  =  13'b1100000011100;     //229pi/512
   cos[229]  =  13'b0000101010001;     //229pi/512
   sin[230]  =  13'b1100000011010;     //230pi/512
   cos[230]  =  13'b0000101000101;     //230pi/512
   sin[231]  =  13'b1100000011000;     //231pi/512
   cos[231]  =  13'b0000100111000;     //231pi/512
   sin[232]  =  13'b1100000010110;     //232pi/512
   cos[232]  =  13'b0000100101100;     //232pi/512
   sin[233]  =  13'b1100000010100;     //233pi/512
   cos[233]  =  13'b0000100100000;     //233pi/512
   sin[234]  =  13'b1100000010011;     //234pi/512
   cos[234]  =  13'b0000100010011;     //234pi/512
   sin[235]  =  13'b1100000010001;     //235pi/512
   cos[235]  =  13'b0000100000111;     //235pi/512
   sin[236]  =  13'b1100000001111;     //236pi/512
   cos[236]  =  13'b0000011111010;     //236pi/512
   sin[237]  =  13'b1100000001110;     //237pi/512
   cos[237]  =  13'b0000011101110;     //237pi/512
   sin[238]  =  13'b1100000001100;     //238pi/512
   cos[238]  =  13'b0000011100001;     //238pi/512
   sin[239]  =  13'b1100000001011;     //239pi/512
   cos[239]  =  13'b0000011010101;     //239pi/512
   sin[240]  =  13'b1100000001010;     //240pi/512
   cos[240]  =  13'b0000011001000;     //240pi/512
   sin[241]  =  13'b1100000001001;     //241pi/512
   cos[241]  =  13'b0000010111100;     //241pi/512
   sin[242]  =  13'b1100000001000;     //242pi/512
   cos[242]  =  13'b0000010101111;     //242pi/512
   sin[243]  =  13'b1100000000111;     //243pi/512
   cos[243]  =  13'b0000010100011;     //243pi/512
   sin[244]  =  13'b1100000000110;     //244pi/512
   cos[244]  =  13'b0000010010110;     //244pi/512
   sin[245]  =  13'b1100000000101;     //245pi/512
   cos[245]  =  13'b0000010001010;     //245pi/512
   sin[246]  =  13'b1100000000100;     //246pi/512
   cos[246]  =  13'b0000001111101;     //246pi/512
   sin[247]  =  13'b1100000000011;     //247pi/512
   cos[247]  =  13'b0000001110001;     //247pi/512
   sin[248]  =  13'b1100000000010;     //248pi/512
   cos[248]  =  13'b0000001100100;     //248pi/512
   sin[249]  =  13'b1100000000010;     //249pi/512
   cos[249]  =  13'b0000001010111;     //249pi/512
   sin[250]  =  13'b1100000000001;     //250pi/512
   cos[250]  =  13'b0000001001011;     //250pi/512
   sin[251]  =  13'b1100000000001;     //251pi/512
   cos[251]  =  13'b0000000111110;     //251pi/512
   sin[252]  =  13'b1100000000001;     //252pi/512
   cos[252]  =  13'b0000000110010;     //252pi/512
   sin[253]  =  13'b1100000000000;     //253pi/512
   cos[253]  =  13'b0000000100101;     //253pi/512
   sin[254]  =  13'b1100000000000;     //254pi/512
   cos[254]  =  13'b0000000011001;     //254pi/512
   sin[255]  =  13'b1100000000000;     //255pi/512
   cos[255]  =  13'b0000000001100;     //255pi/512
   sin[256]  =  13'b1100000000000;     //256pi/512
   cos[256]  =  13'b0000000000000;     //256pi/512
   sin[257]  =  13'b1100000000000;     //257pi/512
   cos[257]  =  13'b1111111110011;     //257pi/512
   sin[258]  =  13'b1100000000000;     //258pi/512
   cos[258]  =  13'b1111111100111;     //258pi/512
   sin[259]  =  13'b1100000000000;     //259pi/512
   cos[259]  =  13'b1111111011010;     //259pi/512
   sin[260]  =  13'b1100000000001;     //260pi/512
   cos[260]  =  13'b1111111001110;     //260pi/512
   sin[261]  =  13'b1100000000001;     //261pi/512
   cos[261]  =  13'b1111111000001;     //261pi/512
   sin[262]  =  13'b1100000000001;     //262pi/512
   cos[262]  =  13'b1111110110101;     //262pi/512
   sin[263]  =  13'b1100000000010;     //263pi/512
   cos[263]  =  13'b1111110101000;     //263pi/512
   sin[264]  =  13'b1100000000010;     //264pi/512
   cos[264]  =  13'b1111110011100;     //264pi/512
   sin[265]  =  13'b1100000000011;     //265pi/512
   cos[265]  =  13'b1111110001111;     //265pi/512
   sin[266]  =  13'b1100000000100;     //266pi/512
   cos[266]  =  13'b1111110000010;     //266pi/512
   sin[267]  =  13'b1100000000101;     //267pi/512
   cos[267]  =  13'b1111101110110;     //267pi/512
   sin[268]  =  13'b1100000000110;     //268pi/512
   cos[268]  =  13'b1111101101001;     //268pi/512
   sin[269]  =  13'b1100000000111;     //269pi/512
   cos[269]  =  13'b1111101011101;     //269pi/512
   sin[270]  =  13'b1100000001000;     //270pi/512
   cos[270]  =  13'b1111101010000;     //270pi/512
   sin[271]  =  13'b1100000001001;     //271pi/512
   cos[271]  =  13'b1111101000100;     //271pi/512
   sin[272]  =  13'b1100000001010;     //272pi/512
   cos[272]  =  13'b1111100110111;     //272pi/512
   sin[273]  =  13'b1100000001011;     //273pi/512
   cos[273]  =  13'b1111100101011;     //273pi/512
   sin[274]  =  13'b1100000001100;     //274pi/512
   cos[274]  =  13'b1111100011110;     //274pi/512
   sin[275]  =  13'b1100000001110;     //275pi/512
   cos[275]  =  13'b1111100010010;     //275pi/512
   sin[276]  =  13'b1100000001111;     //276pi/512
   cos[276]  =  13'b1111100000101;     //276pi/512
   sin[277]  =  13'b1100000010001;     //277pi/512
   cos[277]  =  13'b1111011111001;     //277pi/512
   sin[278]  =  13'b1100000010011;     //278pi/512
   cos[278]  =  13'b1111011101100;     //278pi/512
   sin[279]  =  13'b1100000010100;     //279pi/512
   cos[279]  =  13'b1111011100000;     //279pi/512
   sin[280]  =  13'b1100000010110;     //280pi/512
   cos[280]  =  13'b1111011010011;     //280pi/512
   sin[281]  =  13'b1100000011000;     //281pi/512
   cos[281]  =  13'b1111011000111;     //281pi/512
   sin[282]  =  13'b1100000011010;     //282pi/512
   cos[282]  =  13'b1111010111011;     //282pi/512
   sin[283]  =  13'b1100000011100;     //283pi/512
   cos[283]  =  13'b1111010101110;     //283pi/512
   sin[284]  =  13'b1100000011110;     //284pi/512
   cos[284]  =  13'b1111010100010;     //284pi/512
   sin[285]  =  13'b1100000100000;     //285pi/512
   cos[285]  =  13'b1111010010101;     //285pi/512
   sin[286]  =  13'b1100000100011;     //286pi/512
   cos[286]  =  13'b1111010001001;     //286pi/512
   sin[287]  =  13'b1100000100101;     //287pi/512
   cos[287]  =  13'b1111001111101;     //287pi/512
   sin[288]  =  13'b1100000100111;     //288pi/512
   cos[288]  =  13'b1111001110000;     //288pi/512
   sin[289]  =  13'b1100000101010;     //289pi/512
   cos[289]  =  13'b1111001100100;     //289pi/512
   sin[290]  =  13'b1100000101100;     //290pi/512
   cos[290]  =  13'b1111001011000;     //290pi/512
   sin[291]  =  13'b1100000101111;     //291pi/512
   cos[291]  =  13'b1111001001100;     //291pi/512
   sin[292]  =  13'b1100000110010;     //292pi/512
   cos[292]  =  13'b1111000111111;     //292pi/512
   sin[293]  =  13'b1100000110101;     //293pi/512
   cos[293]  =  13'b1111000110011;     //293pi/512
   sin[294]  =  13'b1100000110111;     //294pi/512
   cos[294]  =  13'b1111000100111;     //294pi/512
   sin[295]  =  13'b1100000111010;     //295pi/512
   cos[295]  =  13'b1111000011011;     //295pi/512
   sin[296]  =  13'b1100000111101;     //296pi/512
   cos[296]  =  13'b1111000001110;     //296pi/512
   sin[297]  =  13'b1100001000000;     //297pi/512
   cos[297]  =  13'b1111000000010;     //297pi/512
   sin[298]  =  13'b1100001000100;     //298pi/512
   cos[298]  =  13'b1110111110110;     //298pi/512
   sin[299]  =  13'b1100001000111;     //299pi/512
   cos[299]  =  13'b1110111101010;     //299pi/512
   sin[300]  =  13'b1100001001010;     //300pi/512
   cos[300]  =  13'b1110111011110;     //300pi/512
   sin[301]  =  13'b1100001001110;     //301pi/512
   cos[301]  =  13'b1110111010010;     //301pi/512
   sin[302]  =  13'b1100001010001;     //302pi/512
   cos[302]  =  13'b1110111000110;     //302pi/512
   sin[303]  =  13'b1100001010101;     //303pi/512
   cos[303]  =  13'b1110110111010;     //303pi/512
   sin[304]  =  13'b1100001011000;     //304pi/512
   cos[304]  =  13'b1110110101101;     //304pi/512
   sin[305]  =  13'b1100001011100;     //305pi/512
   cos[305]  =  13'b1110110100001;     //305pi/512
   sin[306]  =  13'b1100001100000;     //306pi/512
   cos[306]  =  13'b1110110010101;     //306pi/512
   sin[307]  =  13'b1100001100011;     //307pi/512
   cos[307]  =  13'b1110110001010;     //307pi/512
   sin[308]  =  13'b1100001100111;     //308pi/512
   cos[308]  =  13'b1110101111110;     //308pi/512
   sin[309]  =  13'b1100001101011;     //309pi/512
   cos[309]  =  13'b1110101110010;     //309pi/512
   sin[310]  =  13'b1100001101111;     //310pi/512
   cos[310]  =  13'b1110101100110;     //310pi/512
   sin[311]  =  13'b1100001110100;     //311pi/512
   cos[311]  =  13'b1110101011010;     //311pi/512
   sin[312]  =  13'b1100001111000;     //312pi/512
   cos[312]  =  13'b1110101001110;     //312pi/512
   sin[313]  =  13'b1100001111100;     //313pi/512
   cos[313]  =  13'b1110101000010;     //313pi/512
   sin[314]  =  13'b1100010000000;     //314pi/512
   cos[314]  =  13'b1110100110110;     //314pi/512
   sin[315]  =  13'b1100010000101;     //315pi/512
   cos[315]  =  13'b1110100101011;     //315pi/512
   sin[316]  =  13'b1100010001001;     //316pi/512
   cos[316]  =  13'b1110100011111;     //316pi/512
   sin[317]  =  13'b1100010001110;     //317pi/512
   cos[317]  =  13'b1110100010011;     //317pi/512
   sin[318]  =  13'b1100010010010;     //318pi/512
   cos[318]  =  13'b1110100001000;     //318pi/512
   sin[319]  =  13'b1100010010111;     //319pi/512
   cos[319]  =  13'b1110011111100;     //319pi/512
   sin[320]  =  13'b1100010011100;     //320pi/512
   cos[320]  =  13'b1110011110000;     //320pi/512
   sin[321]  =  13'b1100010100001;     //321pi/512
   cos[321]  =  13'b1110011100101;     //321pi/512
   sin[322]  =  13'b1100010100110;     //322pi/512
   cos[322]  =  13'b1110011011001;     //322pi/512
   sin[323]  =  13'b1100010101011;     //323pi/512
   cos[323]  =  13'b1110011001110;     //323pi/512
   sin[324]  =  13'b1100010110000;     //324pi/512
   cos[324]  =  13'b1110011000010;     //324pi/512
   sin[325]  =  13'b1100010110101;     //325pi/512
   cos[325]  =  13'b1110010110111;     //325pi/512
   sin[326]  =  13'b1100010111010;     //326pi/512
   cos[326]  =  13'b1110010101011;     //326pi/512
   sin[327]  =  13'b1100010111111;     //327pi/512
   cos[327]  =  13'b1110010100000;     //327pi/512
   sin[328]  =  13'b1100011000101;     //328pi/512
   cos[328]  =  13'b1110010010100;     //328pi/512
   sin[329]  =  13'b1100011001010;     //329pi/512
   cos[329]  =  13'b1110010001001;     //329pi/512
   sin[330]  =  13'b1100011010000;     //330pi/512
   cos[330]  =  13'b1110001111110;     //330pi/512
   sin[331]  =  13'b1100011010101;     //331pi/512
   cos[331]  =  13'b1110001110010;     //331pi/512
   sin[332]  =  13'b1100011011011;     //332pi/512
   cos[332]  =  13'b1110001100111;     //332pi/512
   sin[333]  =  13'b1100011100000;     //333pi/512
   cos[333]  =  13'b1110001011100;     //333pi/512
   sin[334]  =  13'b1100011100110;     //334pi/512
   cos[334]  =  13'b1110001010001;     //334pi/512
   sin[335]  =  13'b1100011101100;     //335pi/512
   cos[335]  =  13'b1110001000110;     //335pi/512
   sin[336]  =  13'b1100011110010;     //336pi/512
   cos[336]  =  13'b1110000111011;     //336pi/512
   sin[337]  =  13'b1100011111000;     //337pi/512
   cos[337]  =  13'b1110000110000;     //337pi/512
   sin[338]  =  13'b1100011111110;     //338pi/512
   cos[338]  =  13'b1110000100100;     //338pi/512
   sin[339]  =  13'b1100100000100;     //339pi/512
   cos[339]  =  13'b1110000011001;     //339pi/512
   sin[340]  =  13'b1100100001010;     //340pi/512
   cos[340]  =  13'b1110000001111;     //340pi/512
   sin[341]  =  13'b1100100010000;     //341pi/512
   cos[341]  =  13'b1110000000100;     //341pi/512
   sin[342]  =  13'b1100100010111;     //342pi/512
   cos[342]  =  13'b1101111111001;     //342pi/512
   sin[343]  =  13'b1100100011101;     //343pi/512
   cos[343]  =  13'b1101111101110;     //343pi/512
   sin[344]  =  13'b1100100100011;     //344pi/512
   cos[344]  =  13'b1101111100011;     //344pi/512
   sin[345]  =  13'b1100100101010;     //345pi/512
   cos[345]  =  13'b1101111011000;     //345pi/512
   sin[346]  =  13'b1100100110000;     //346pi/512
   cos[346]  =  13'b1101111001110;     //346pi/512
   sin[347]  =  13'b1100100110111;     //347pi/512
   cos[347]  =  13'b1101111000011;     //347pi/512
   sin[348]  =  13'b1100100111110;     //348pi/512
   cos[348]  =  13'b1101110111000;     //348pi/512
   sin[349]  =  13'b1100101000100;     //349pi/512
   cos[349]  =  13'b1101110101110;     //349pi/512
   sin[350]  =  13'b1100101001011;     //350pi/512
   cos[350]  =  13'b1101110100011;     //350pi/512
   sin[351]  =  13'b1100101010010;     //351pi/512
   cos[351]  =  13'b1101110011001;     //351pi/512
   sin[352]  =  13'b1100101011001;     //352pi/512
   cos[352]  =  13'b1101110001110;     //352pi/512
   sin[353]  =  13'b1100101100000;     //353pi/512
   cos[353]  =  13'b1101110000100;     //353pi/512
   sin[354]  =  13'b1100101100111;     //354pi/512
   cos[354]  =  13'b1101101111001;     //354pi/512
   sin[355]  =  13'b1100101101110;     //355pi/512
   cos[355]  =  13'b1101101101111;     //355pi/512
   sin[356]  =  13'b1100101110110;     //356pi/512
   cos[356]  =  13'b1101101100101;     //356pi/512
   sin[357]  =  13'b1100101111101;     //357pi/512
   cos[357]  =  13'b1101101011010;     //357pi/512
   sin[358]  =  13'b1100110000100;     //358pi/512
   cos[358]  =  13'b1101101010000;     //358pi/512
   sin[359]  =  13'b1100110001100;     //359pi/512
   cos[359]  =  13'b1101101000110;     //359pi/512
   sin[360]  =  13'b1100110010011;     //360pi/512
   cos[360]  =  13'b1101100111100;     //360pi/512
   sin[361]  =  13'b1100110011011;     //361pi/512
   cos[361]  =  13'b1101100110010;     //361pi/512
   sin[362]  =  13'b1100110100010;     //362pi/512
   cos[362]  =  13'b1101100101000;     //362pi/512
   sin[363]  =  13'b1100110101010;     //363pi/512
   cos[363]  =  13'b1101100011110;     //363pi/512
   sin[364]  =  13'b1100110110001;     //364pi/512
   cos[364]  =  13'b1101100010100;     //364pi/512
   sin[365]  =  13'b1100110111001;     //365pi/512
   cos[365]  =  13'b1101100001010;     //365pi/512
   sin[366]  =  13'b1100111000001;     //366pi/512
   cos[366]  =  13'b1101100000000;     //366pi/512
   sin[367]  =  13'b1100111001001;     //367pi/512
   cos[367]  =  13'b1101011110111;     //367pi/512
   sin[368]  =  13'b1100111010001;     //368pi/512
   cos[368]  =  13'b1101011101101;     //368pi/512
   sin[369]  =  13'b1100111011001;     //369pi/512
   cos[369]  =  13'b1101011100011;     //369pi/512
   sin[370]  =  13'b1100111100001;     //370pi/512
   cos[370]  =  13'b1101011011001;     //370pi/512
   sin[371]  =  13'b1100111101001;     //371pi/512
   cos[371]  =  13'b1101011010000;     //371pi/512
   sin[372]  =  13'b1100111110001;     //372pi/512
   cos[372]  =  13'b1101011000110;     //372pi/512
   sin[373]  =  13'b1100111111001;     //373pi/512
   cos[373]  =  13'b1101010111101;     //373pi/512
   sin[374]  =  13'b1101000000010;     //374pi/512
   cos[374]  =  13'b1101010110011;     //374pi/512
   sin[375]  =  13'b1101000001010;     //375pi/512
   cos[375]  =  13'b1101010101010;     //375pi/512
   sin[376]  =  13'b1101000010011;     //376pi/512
   cos[376]  =  13'b1101010100001;     //376pi/512
   sin[377]  =  13'b1101000011011;     //377pi/512
   cos[377]  =  13'b1101010010111;     //377pi/512
   sin[378]  =  13'b1101000100100;     //378pi/512
   cos[378]  =  13'b1101010001110;     //378pi/512
   sin[379]  =  13'b1101000101100;     //379pi/512
   cos[379]  =  13'b1101010000101;     //379pi/512
   sin[380]  =  13'b1101000110101;     //380pi/512
   cos[380]  =  13'b1101001111100;     //380pi/512
   sin[381]  =  13'b1101000111101;     //381pi/512
   cos[381]  =  13'b1101001110011;     //381pi/512
   sin[382]  =  13'b1101001000110;     //382pi/512
   cos[382]  =  13'b1101001101010;     //382pi/512
   sin[383]  =  13'b1101001001111;     //383pi/512
   cos[383]  =  13'b1101001100001;     //383pi/512
   sin[384]  =  13'b1101001011000;     //384pi/512
   cos[384]  =  13'b1101001011000;     //384pi/512
   sin[385]  =  13'b1101001100001;     //385pi/512
   cos[385]  =  13'b1101001001111;     //385pi/512
   sin[386]  =  13'b1101001101010;     //386pi/512
   cos[386]  =  13'b1101001000110;     //386pi/512
   sin[387]  =  13'b1101001110011;     //387pi/512
   cos[387]  =  13'b1101000111101;     //387pi/512
   sin[388]  =  13'b1101001111100;     //388pi/512
   cos[388]  =  13'b1101000110101;     //388pi/512
   sin[389]  =  13'b1101010000101;     //389pi/512
   cos[389]  =  13'b1101000101100;     //389pi/512
   sin[390]  =  13'b1101010001110;     //390pi/512
   cos[390]  =  13'b1101000100100;     //390pi/512
   sin[391]  =  13'b1101010010111;     //391pi/512
   cos[391]  =  13'b1101000011011;     //391pi/512
   sin[392]  =  13'b1101010100001;     //392pi/512
   cos[392]  =  13'b1101000010011;     //392pi/512
   sin[393]  =  13'b1101010101010;     //393pi/512
   cos[393]  =  13'b1101000001010;     //393pi/512
   sin[394]  =  13'b1101010110011;     //394pi/512
   cos[394]  =  13'b1101000000010;     //394pi/512
   sin[395]  =  13'b1101010111101;     //395pi/512
   cos[395]  =  13'b1100111111001;     //395pi/512
   sin[396]  =  13'b1101011000110;     //396pi/512
   cos[396]  =  13'b1100111110001;     //396pi/512
   sin[397]  =  13'b1101011010000;     //397pi/512
   cos[397]  =  13'b1100111101001;     //397pi/512
   sin[398]  =  13'b1101011011001;     //398pi/512
   cos[398]  =  13'b1100111100001;     //398pi/512
   sin[399]  =  13'b1101011100011;     //399pi/512
   cos[399]  =  13'b1100111011001;     //399pi/512
   sin[400]  =  13'b1101011101101;     //400pi/512
   cos[400]  =  13'b1100111010001;     //400pi/512
   sin[401]  =  13'b1101011110111;     //401pi/512
   cos[401]  =  13'b1100111001001;     //401pi/512
   sin[402]  =  13'b1101100000000;     //402pi/512
   cos[402]  =  13'b1100111000001;     //402pi/512
   sin[403]  =  13'b1101100001010;     //403pi/512
   cos[403]  =  13'b1100110111001;     //403pi/512
   sin[404]  =  13'b1101100010100;     //404pi/512
   cos[404]  =  13'b1100110110001;     //404pi/512
   sin[405]  =  13'b1101100011110;     //405pi/512
   cos[405]  =  13'b1100110101010;     //405pi/512
   sin[406]  =  13'b1101100101000;     //406pi/512
   cos[406]  =  13'b1100110100010;     //406pi/512
   sin[407]  =  13'b1101100110010;     //407pi/512
   cos[407]  =  13'b1100110011011;     //407pi/512
   sin[408]  =  13'b1101100111100;     //408pi/512
   cos[408]  =  13'b1100110010011;     //408pi/512
   sin[409]  =  13'b1101101000110;     //409pi/512
   cos[409]  =  13'b1100110001100;     //409pi/512
   sin[410]  =  13'b1101101010000;     //410pi/512
   cos[410]  =  13'b1100110000100;     //410pi/512
   sin[411]  =  13'b1101101011010;     //411pi/512
   cos[411]  =  13'b1100101111101;     //411pi/512
   sin[412]  =  13'b1101101100101;     //412pi/512
   cos[412]  =  13'b1100101110110;     //412pi/512
   sin[413]  =  13'b1101101101111;     //413pi/512
   cos[413]  =  13'b1100101101110;     //413pi/512
   sin[414]  =  13'b1101101111001;     //414pi/512
   cos[414]  =  13'b1100101100111;     //414pi/512
   sin[415]  =  13'b1101110000100;     //415pi/512
   cos[415]  =  13'b1100101100000;     //415pi/512
   sin[416]  =  13'b1101110001110;     //416pi/512
   cos[416]  =  13'b1100101011001;     //416pi/512
   sin[417]  =  13'b1101110011001;     //417pi/512
   cos[417]  =  13'b1100101010010;     //417pi/512
   sin[418]  =  13'b1101110100011;     //418pi/512
   cos[418]  =  13'b1100101001011;     //418pi/512
   sin[419]  =  13'b1101110101110;     //419pi/512
   cos[419]  =  13'b1100101000100;     //419pi/512
   sin[420]  =  13'b1101110111000;     //420pi/512
   cos[420]  =  13'b1100100111110;     //420pi/512
   sin[421]  =  13'b1101111000011;     //421pi/512
   cos[421]  =  13'b1100100110111;     //421pi/512
   sin[422]  =  13'b1101111001110;     //422pi/512
   cos[422]  =  13'b1100100110000;     //422pi/512
   sin[423]  =  13'b1101111011000;     //423pi/512
   cos[423]  =  13'b1100100101010;     //423pi/512
   sin[424]  =  13'b1101111100011;     //424pi/512
   cos[424]  =  13'b1100100100011;     //424pi/512
   sin[425]  =  13'b1101111101110;     //425pi/512
   cos[425]  =  13'b1100100011101;     //425pi/512
   sin[426]  =  13'b1101111111001;     //426pi/512
   cos[426]  =  13'b1100100010111;     //426pi/512
   sin[427]  =  13'b1110000000100;     //427pi/512
   cos[427]  =  13'b1100100010000;     //427pi/512
   sin[428]  =  13'b1110000001111;     //428pi/512
   cos[428]  =  13'b1100100001010;     //428pi/512
   sin[429]  =  13'b1110000011001;     //429pi/512
   cos[429]  =  13'b1100100000100;     //429pi/512
   sin[430]  =  13'b1110000100100;     //430pi/512
   cos[430]  =  13'b1100011111110;     //430pi/512
   sin[431]  =  13'b1110000110000;     //431pi/512
   cos[431]  =  13'b1100011111000;     //431pi/512
   sin[432]  =  13'b1110000111011;     //432pi/512
   cos[432]  =  13'b1100011110010;     //432pi/512
   sin[433]  =  13'b1110001000110;     //433pi/512
   cos[433]  =  13'b1100011101100;     //433pi/512
   sin[434]  =  13'b1110001010001;     //434pi/512
   cos[434]  =  13'b1100011100110;     //434pi/512
   sin[435]  =  13'b1110001011100;     //435pi/512
   cos[435]  =  13'b1100011100000;     //435pi/512
   sin[436]  =  13'b1110001100111;     //436pi/512
   cos[436]  =  13'b1100011011011;     //436pi/512
   sin[437]  =  13'b1110001110010;     //437pi/512
   cos[437]  =  13'b1100011010101;     //437pi/512
   sin[438]  =  13'b1110001111110;     //438pi/512
   cos[438]  =  13'b1100011010000;     //438pi/512
   sin[439]  =  13'b1110010001001;     //439pi/512
   cos[439]  =  13'b1100011001010;     //439pi/512
   sin[440]  =  13'b1110010010100;     //440pi/512
   cos[440]  =  13'b1100011000101;     //440pi/512
   sin[441]  =  13'b1110010100000;     //441pi/512
   cos[441]  =  13'b1100010111111;     //441pi/512
   sin[442]  =  13'b1110010101011;     //442pi/512
   cos[442]  =  13'b1100010111010;     //442pi/512
   sin[443]  =  13'b1110010110111;     //443pi/512
   cos[443]  =  13'b1100010110101;     //443pi/512
   sin[444]  =  13'b1110011000010;     //444pi/512
   cos[444]  =  13'b1100010110000;     //444pi/512
   sin[445]  =  13'b1110011001110;     //445pi/512
   cos[445]  =  13'b1100010101011;     //445pi/512
   sin[446]  =  13'b1110011011001;     //446pi/512
   cos[446]  =  13'b1100010100110;     //446pi/512
   sin[447]  =  13'b1110011100101;     //447pi/512
   cos[447]  =  13'b1100010100001;     //447pi/512
   sin[448]  =  13'b1110011110000;     //448pi/512
   cos[448]  =  13'b1100010011100;     //448pi/512
   sin[449]  =  13'b1110011111100;     //449pi/512
   cos[449]  =  13'b1100010010111;     //449pi/512
   sin[450]  =  13'b1110100001000;     //450pi/512
   cos[450]  =  13'b1100010010010;     //450pi/512
   sin[451]  =  13'b1110100010011;     //451pi/512
   cos[451]  =  13'b1100010001110;     //451pi/512
   sin[452]  =  13'b1110100011111;     //452pi/512
   cos[452]  =  13'b1100010001001;     //452pi/512
   sin[453]  =  13'b1110100101011;     //453pi/512
   cos[453]  =  13'b1100010000101;     //453pi/512
   sin[454]  =  13'b1110100110110;     //454pi/512
   cos[454]  =  13'b1100010000000;     //454pi/512
   sin[455]  =  13'b1110101000010;     //455pi/512
   cos[455]  =  13'b1100001111100;     //455pi/512
   sin[456]  =  13'b1110101001110;     //456pi/512
   cos[456]  =  13'b1100001111000;     //456pi/512
   sin[457]  =  13'b1110101011010;     //457pi/512
   cos[457]  =  13'b1100001110100;     //457pi/512
   sin[458]  =  13'b1110101100110;     //458pi/512
   cos[458]  =  13'b1100001101111;     //458pi/512
   sin[459]  =  13'b1110101110010;     //459pi/512
   cos[459]  =  13'b1100001101011;     //459pi/512
   sin[460]  =  13'b1110101111110;     //460pi/512
   cos[460]  =  13'b1100001100111;     //460pi/512
   sin[461]  =  13'b1110110001010;     //461pi/512
   cos[461]  =  13'b1100001100011;     //461pi/512
   sin[462]  =  13'b1110110010101;     //462pi/512
   cos[462]  =  13'b1100001100000;     //462pi/512
   sin[463]  =  13'b1110110100001;     //463pi/512
   cos[463]  =  13'b1100001011100;     //463pi/512
   sin[464]  =  13'b1110110101101;     //464pi/512
   cos[464]  =  13'b1100001011000;     //464pi/512
   sin[465]  =  13'b1110110111010;     //465pi/512
   cos[465]  =  13'b1100001010101;     //465pi/512
   sin[466]  =  13'b1110111000110;     //466pi/512
   cos[466]  =  13'b1100001010001;     //466pi/512
   sin[467]  =  13'b1110111010010;     //467pi/512
   cos[467]  =  13'b1100001001110;     //467pi/512
   sin[468]  =  13'b1110111011110;     //468pi/512
   cos[468]  =  13'b1100001001010;     //468pi/512
   sin[469]  =  13'b1110111101010;     //469pi/512
   cos[469]  =  13'b1100001000111;     //469pi/512
   sin[470]  =  13'b1110111110110;     //470pi/512
   cos[470]  =  13'b1100001000100;     //470pi/512
   sin[471]  =  13'b1111000000010;     //471pi/512
   cos[471]  =  13'b1100001000000;     //471pi/512
   sin[472]  =  13'b1111000001110;     //472pi/512
   cos[472]  =  13'b1100000111101;     //472pi/512
   sin[473]  =  13'b1111000011011;     //473pi/512
   cos[473]  =  13'b1100000111010;     //473pi/512
   sin[474]  =  13'b1111000100111;     //474pi/512
   cos[474]  =  13'b1100000110111;     //474pi/512
   sin[475]  =  13'b1111000110011;     //475pi/512
   cos[475]  =  13'b1100000110101;     //475pi/512
   sin[476]  =  13'b1111000111111;     //476pi/512
   cos[476]  =  13'b1100000110010;     //476pi/512
   sin[477]  =  13'b1111001001100;     //477pi/512
   cos[477]  =  13'b1100000101111;     //477pi/512
   sin[478]  =  13'b1111001011000;     //478pi/512
   cos[478]  =  13'b1100000101100;     //478pi/512
   sin[479]  =  13'b1111001100100;     //479pi/512
   cos[479]  =  13'b1100000101010;     //479pi/512
   sin[480]  =  13'b1111001110000;     //480pi/512
   cos[480]  =  13'b1100000100111;     //480pi/512
   sin[481]  =  13'b1111001111101;     //481pi/512
   cos[481]  =  13'b1100000100101;     //481pi/512
   sin[482]  =  13'b1111010001001;     //482pi/512
   cos[482]  =  13'b1100000100011;     //482pi/512
   sin[483]  =  13'b1111010010101;     //483pi/512
   cos[483]  =  13'b1100000100000;     //483pi/512
   sin[484]  =  13'b1111010100010;     //484pi/512
   cos[484]  =  13'b1100000011110;     //484pi/512
   sin[485]  =  13'b1111010101110;     //485pi/512
   cos[485]  =  13'b1100000011100;     //485pi/512
   sin[486]  =  13'b1111010111011;     //486pi/512
   cos[486]  =  13'b1100000011010;     //486pi/512
   sin[487]  =  13'b1111011000111;     //487pi/512
   cos[487]  =  13'b1100000011000;     //487pi/512
   sin[488]  =  13'b1111011010011;     //488pi/512
   cos[488]  =  13'b1100000010110;     //488pi/512
   sin[489]  =  13'b1111011100000;     //489pi/512
   cos[489]  =  13'b1100000010100;     //489pi/512
   sin[490]  =  13'b1111011101100;     //490pi/512
   cos[490]  =  13'b1100000010011;     //490pi/512
   sin[491]  =  13'b1111011111001;     //491pi/512
   cos[491]  =  13'b1100000010001;     //491pi/512
   sin[492]  =  13'b1111100000101;     //492pi/512
   cos[492]  =  13'b1100000001111;     //492pi/512
   sin[493]  =  13'b1111100010010;     //493pi/512
   cos[493]  =  13'b1100000001110;     //493pi/512
   sin[494]  =  13'b1111100011110;     //494pi/512
   cos[494]  =  13'b1100000001100;     //494pi/512
   sin[495]  =  13'b1111100101011;     //495pi/512
   cos[495]  =  13'b1100000001011;     //495pi/512
   sin[496]  =  13'b1111100110111;     //496pi/512
   cos[496]  =  13'b1100000001010;     //496pi/512
   sin[497]  =  13'b1111101000100;     //497pi/512
   cos[497]  =  13'b1100000001001;     //497pi/512
   sin[498]  =  13'b1111101010000;     //498pi/512
   cos[498]  =  13'b1100000001000;     //498pi/512
   sin[499]  =  13'b1111101011101;     //499pi/512
   cos[499]  =  13'b1100000000111;     //499pi/512
   sin[500]  =  13'b1111101101001;     //500pi/512
   cos[500]  =  13'b1100000000110;     //500pi/512
   sin[501]  =  13'b1111101110110;     //501pi/512
   cos[501]  =  13'b1100000000101;     //501pi/512
   sin[502]  =  13'b1111110000010;     //502pi/512
   cos[502]  =  13'b1100000000100;     //502pi/512
   sin[503]  =  13'b1111110001111;     //503pi/512
   cos[503]  =  13'b1100000000011;     //503pi/512
   sin[504]  =  13'b1111110011100;     //504pi/512
   cos[504]  =  13'b1100000000010;     //504pi/512
   sin[505]  =  13'b1111110101000;     //505pi/512
   cos[505]  =  13'b1100000000010;     //505pi/512
   sin[506]  =  13'b1111110110101;     //506pi/512
   cos[506]  =  13'b1100000000001;     //506pi/512
   sin[507]  =  13'b1111111000001;     //507pi/512
   cos[507]  =  13'b1100000000001;     //507pi/512
   sin[508]  =  13'b1111111001110;     //508pi/512
   cos[508]  =  13'b1100000000001;     //508pi/512
   sin[509]  =  13'b1111111011010;     //509pi/512
   cos[509]  =  13'b1100000000000;     //509pi/512
   sin[510]  =  13'b1111111100111;     //510pi/512
   cos[510]  =  13'b1100000000000;     //510pi/512
   sin[511]  =  13'b1111111110011;     //511pi/512
   cos[511]  =  13'b1100000000000;     //511pi/512
   m_sin[0]  =  13'b0000000000000;     //0pi/512
   m_cos[0]  =  13'b0100000000000;     //0pi/512
   m_sin[1]  =  13'b1111111110101;     //1pi/512
   m_cos[1]  =  13'b0011111111111;     //1pi/512
   m_sin[2]  =  13'b1111111101001;     //2pi/512
   m_cos[2]  =  13'b0011111111111;     //2pi/512
   m_sin[3]  =  13'b1111111011110;     //3pi/512
   m_cos[3]  =  13'b0011111111111;     //3pi/512
   m_sin[4]  =  13'b1111111010011;     //4pi/512
   m_cos[4]  =  13'b0011111111111;     //4pi/512
   m_sin[5]  =  13'b1111111000111;     //5pi/512
   m_cos[5]  =  13'b0011111111111;     //5pi/512
   m_sin[6]  =  13'b1111110111100;     //6pi/512
   m_cos[6]  =  13'b0011111111110;     //6pi/512
   m_sin[7]  =  13'b1111110110001;     //7pi/512
   m_cos[7]  =  13'b0011111111110;     //7pi/512
   m_sin[8]  =  13'b1111110100110;     //8pi/512
   m_cos[8]  =  13'b0011111111110;     //8pi/512
   m_sin[9]  =  13'b1111110011010;     //9pi/512
   m_cos[9]  =  13'b0011111111101;     //9pi/512
   m_sin[10]  =  13'b1111110001111;     //10pi/512
   m_cos[10]  =  13'b0011111111100;     //10pi/512
   m_sin[11]  =  13'b1111110000100;     //11pi/512
   m_cos[11]  =  13'b0011111111100;     //11pi/512
   m_sin[12]  =  13'b1111101111000;     //12pi/512
   m_cos[12]  =  13'b0011111111011;     //12pi/512
   m_sin[13]  =  13'b1111101101101;     //13pi/512
   m_cos[13]  =  13'b0011111111010;     //13pi/512
   m_sin[14]  =  13'b1111101100010;     //14pi/512
   m_cos[14]  =  13'b0011111111001;     //14pi/512
   m_sin[15]  =  13'b1111101010111;     //15pi/512
   m_cos[15]  =  13'b0011111111000;     //15pi/512
   m_sin[16]  =  13'b1111101001011;     //16pi/512
   m_cos[16]  =  13'b0011111111000;     //16pi/512
   m_sin[17]  =  13'b1111101000000;     //17pi/512
   m_cos[17]  =  13'b0011111110110;     //17pi/512
   m_sin[18]  =  13'b1111100110101;     //18pi/512
   m_cos[18]  =  13'b0011111110101;     //18pi/512
   m_sin[19]  =  13'b1111100101010;     //19pi/512
   m_cos[19]  =  13'b0011111110100;     //19pi/512
   m_sin[20]  =  13'b1111100011110;     //20pi/512
   m_cos[20]  =  13'b0011111110011;     //20pi/512
   m_sin[21]  =  13'b1111100010011;     //21pi/512
   m_cos[21]  =  13'b0011111110010;     //21pi/512
   m_sin[22]  =  13'b1111100001000;     //22pi/512
   m_cos[22]  =  13'b0011111110000;     //22pi/512
   m_sin[23]  =  13'b1111011111101;     //23pi/512
   m_cos[23]  =  13'b0011111101111;     //23pi/512
   m_sin[24]  =  13'b1111011110001;     //24pi/512
   m_cos[24]  =  13'b0011111101110;     //24pi/512
   m_sin[25]  =  13'b1111011100110;     //25pi/512
   m_cos[25]  =  13'b0011111101100;     //25pi/512
   m_sin[26]  =  13'b1111011011011;     //26pi/512
   m_cos[26]  =  13'b0011111101010;     //26pi/512
   m_sin[27]  =  13'b1111011010000;     //27pi/512
   m_cos[27]  =  13'b0011111101001;     //27pi/512
   m_sin[28]  =  13'b1111011000101;     //28pi/512
   m_cos[28]  =  13'b0011111100111;     //28pi/512
   m_sin[29]  =  13'b1111010111001;     //29pi/512
   m_cos[29]  =  13'b0011111100101;     //29pi/512
   m_sin[30]  =  13'b1111010101110;     //30pi/512
   m_cos[30]  =  13'b0011111100011;     //30pi/512
   m_sin[31]  =  13'b1111010100011;     //31pi/512
   m_cos[31]  =  13'b0011111100010;     //31pi/512
   m_sin[32]  =  13'b1111010011000;     //32pi/512
   m_cos[32]  =  13'b0011111100000;     //32pi/512
   m_sin[33]  =  13'b1111010001101;     //33pi/512
   m_cos[33]  =  13'b0011111011110;     //33pi/512
   m_sin[34]  =  13'b1111010000010;     //34pi/512
   m_cos[34]  =  13'b0011111011100;     //34pi/512
   m_sin[35]  =  13'b1111001110111;     //35pi/512
   m_cos[35]  =  13'b0011111011001;     //35pi/512
   m_sin[36]  =  13'b1111001101100;     //36pi/512
   m_cos[36]  =  13'b0011111010111;     //36pi/512
   m_sin[37]  =  13'b1111001100000;     //37pi/512
   m_cos[37]  =  13'b0011111010101;     //37pi/512
   m_sin[38]  =  13'b1111001010101;     //38pi/512
   m_cos[38]  =  13'b0011111010011;     //38pi/512
   m_sin[39]  =  13'b1111001001010;     //39pi/512
   m_cos[39]  =  13'b0011111010000;     //39pi/512
   m_sin[40]  =  13'b1111000111111;     //40pi/512
   m_cos[40]  =  13'b0011111001110;     //40pi/512
   m_sin[41]  =  13'b1111000110100;     //41pi/512
   m_cos[41]  =  13'b0011111001011;     //41pi/512
   m_sin[42]  =  13'b1111000101001;     //42pi/512
   m_cos[42]  =  13'b0011111001001;     //42pi/512
   m_sin[43]  =  13'b1111000011110;     //43pi/512
   m_cos[43]  =  13'b0011111000110;     //43pi/512
   m_sin[44]  =  13'b1111000010011;     //44pi/512
   m_cos[44]  =  13'b0011111000011;     //44pi/512
   m_sin[45]  =  13'b1111000001000;     //45pi/512
   m_cos[45]  =  13'b0011111000001;     //45pi/512
   m_sin[46]  =  13'b1110111111101;     //46pi/512
   m_cos[46]  =  13'b0011110111110;     //46pi/512
   m_sin[47]  =  13'b1110111110010;     //47pi/512
   m_cos[47]  =  13'b0011110111011;     //47pi/512
   m_sin[48]  =  13'b1110111100111;     //48pi/512
   m_cos[48]  =  13'b0011110111000;     //48pi/512
   m_sin[49]  =  13'b1110111011101;     //49pi/512
   m_cos[49]  =  13'b0011110110101;     //49pi/512
   m_sin[50]  =  13'b1110111010010;     //50pi/512
   m_cos[50]  =  13'b0011110110010;     //50pi/512
   m_sin[51]  =  13'b1110111000111;     //51pi/512
   m_cos[51]  =  13'b0011110101111;     //51pi/512
   m_sin[52]  =  13'b1110110111100;     //52pi/512
   m_cos[52]  =  13'b0011110101100;     //52pi/512
   m_sin[53]  =  13'b1110110110001;     //53pi/512
   m_cos[53]  =  13'b0011110101000;     //53pi/512
   m_sin[54]  =  13'b1110110100110;     //54pi/512
   m_cos[54]  =  13'b0011110100101;     //54pi/512
   m_sin[55]  =  13'b1110110011011;     //55pi/512
   m_cos[55]  =  13'b0011110100010;     //55pi/512
   m_sin[56]  =  13'b1110110010001;     //56pi/512
   m_cos[56]  =  13'b0011110011110;     //56pi/512
   m_sin[57]  =  13'b1110110000110;     //57pi/512
   m_cos[57]  =  13'b0011110011011;     //57pi/512
   m_sin[58]  =  13'b1110101111011;     //58pi/512
   m_cos[58]  =  13'b0011110010111;     //58pi/512
   m_sin[59]  =  13'b1110101110000;     //59pi/512
   m_cos[59]  =  13'b0011110010100;     //59pi/512
   m_sin[60]  =  13'b1110101100110;     //60pi/512
   m_cos[60]  =  13'b0011110010000;     //60pi/512
   m_sin[61]  =  13'b1110101011011;     //61pi/512
   m_cos[61]  =  13'b0011110001100;     //61pi/512
   m_sin[62]  =  13'b1110101010000;     //62pi/512
   m_cos[62]  =  13'b0011110001001;     //62pi/512
   m_sin[63]  =  13'b1110101000110;     //63pi/512
   m_cos[63]  =  13'b0011110000101;     //63pi/512
   m_sin[64]  =  13'b1110100111011;     //64pi/512
   m_cos[64]  =  13'b0011110000001;     //64pi/512
   m_sin[65]  =  13'b1110100110001;     //65pi/512
   m_cos[65]  =  13'b0011101111101;     //65pi/512
   m_sin[66]  =  13'b1110100100110;     //66pi/512
   m_cos[66]  =  13'b0011101111001;     //66pi/512
   m_sin[67]  =  13'b1110100011011;     //67pi/512
   m_cos[67]  =  13'b0011101110101;     //67pi/512
   m_sin[68]  =  13'b1110100010001;     //68pi/512
   m_cos[68]  =  13'b0011101110001;     //68pi/512
   m_sin[69]  =  13'b1110100000110;     //69pi/512
   m_cos[69]  =  13'b0011101101101;     //69pi/512
   m_sin[70]  =  13'b1110011111100;     //70pi/512
   m_cos[70]  =  13'b0011101101000;     //70pi/512
   m_sin[71]  =  13'b1110011110001;     //71pi/512
   m_cos[71]  =  13'b0011101100100;     //71pi/512
   m_sin[72]  =  13'b1110011100111;     //72pi/512
   m_cos[72]  =  13'b0011101100000;     //72pi/512
   m_sin[73]  =  13'b1110011011101;     //73pi/512
   m_cos[73]  =  13'b0011101011011;     //73pi/512
   m_sin[74]  =  13'b1110011010010;     //74pi/512
   m_cos[74]  =  13'b0011101010111;     //74pi/512
   m_sin[75]  =  13'b1110011001000;     //75pi/512
   m_cos[75]  =  13'b0011101010010;     //75pi/512
   m_sin[76]  =  13'b1110010111101;     //76pi/512
   m_cos[76]  =  13'b0011101001110;     //76pi/512
   m_sin[77]  =  13'b1110010110011;     //77pi/512
   m_cos[77]  =  13'b0011101001001;     //77pi/512
   m_sin[78]  =  13'b1110010101001;     //78pi/512
   m_cos[78]  =  13'b0011101000100;     //78pi/512
   m_sin[79]  =  13'b1110010011111;     //79pi/512
   m_cos[79]  =  13'b0011101000000;     //79pi/512
   m_sin[80]  =  13'b1110010010100;     //80pi/512
   m_cos[80]  =  13'b0011100111011;     //80pi/512
   m_sin[81]  =  13'b1110010001010;     //81pi/512
   m_cos[81]  =  13'b0011100110110;     //81pi/512
   m_sin[82]  =  13'b1110010000000;     //82pi/512
   m_cos[82]  =  13'b0011100110001;     //82pi/512
   m_sin[83]  =  13'b1110001110110;     //83pi/512
   m_cos[83]  =  13'b0011100101100;     //83pi/512
   m_sin[84]  =  13'b1110001101100;     //84pi/512
   m_cos[84]  =  13'b0011100100111;     //84pi/512
   m_sin[85]  =  13'b1110001100010;     //85pi/512
   m_cos[85]  =  13'b0011100100010;     //85pi/512
   m_sin[86]  =  13'b1110001011000;     //86pi/512
   m_cos[86]  =  13'b0011100011101;     //86pi/512
   m_sin[87]  =  13'b1110001001101;     //87pi/512
   m_cos[87]  =  13'b0011100011000;     //87pi/512
   m_sin[88]  =  13'b1110001000011;     //88pi/512
   m_cos[88]  =  13'b0011100010010;     //88pi/512
   m_sin[89]  =  13'b1110000111001;     //89pi/512
   m_cos[89]  =  13'b0011100001101;     //89pi/512
   m_sin[90]  =  13'b1110000110000;     //90pi/512
   m_cos[90]  =  13'b0011100001000;     //90pi/512
   m_sin[91]  =  13'b1110000100110;     //91pi/512
   m_cos[91]  =  13'b0011100000010;     //91pi/512
   m_sin[92]  =  13'b1110000011100;     //92pi/512
   m_cos[92]  =  13'b0011011111101;     //92pi/512
   m_sin[93]  =  13'b1110000010010;     //93pi/512
   m_cos[93]  =  13'b0011011110111;     //93pi/512
   m_sin[94]  =  13'b1110000001000;     //94pi/512
   m_cos[94]  =  13'b0011011110010;     //94pi/512
   m_sin[95]  =  13'b1101111111110;     //95pi/512
   m_cos[95]  =  13'b0011011101100;     //95pi/512
   m_sin[96]  =  13'b1101111110100;     //96pi/512
   m_cos[96]  =  13'b0011011100110;     //96pi/512
   m_sin[97]  =  13'b1101111101011;     //97pi/512
   m_cos[97]  =  13'b0011011100001;     //97pi/512
   m_sin[98]  =  13'b1101111100001;     //98pi/512
   m_cos[98]  =  13'b0011011011011;     //98pi/512
   m_sin[99]  =  13'b1101111010111;     //99pi/512
   m_cos[99]  =  13'b0011011010101;     //99pi/512
   m_sin[100]  =  13'b1101111001110;     //100pi/512
   m_cos[100]  =  13'b0011011001111;     //100pi/512
   m_sin[101]  =  13'b1101111000100;     //101pi/512
   m_cos[101]  =  13'b0011011001001;     //101pi/512
   m_sin[102]  =  13'b1101110111010;     //102pi/512
   m_cos[102]  =  13'b0011011000011;     //102pi/512
   m_sin[103]  =  13'b1101110110001;     //103pi/512
   m_cos[103]  =  13'b0011010111101;     //103pi/512
   m_sin[104]  =  13'b1101110100111;     //104pi/512
   m_cos[104]  =  13'b0011010110111;     //104pi/512
   m_sin[105]  =  13'b1101110011110;     //105pi/512
   m_cos[105]  =  13'b0011010110001;     //105pi/512
   m_sin[106]  =  13'b1101110010100;     //106pi/512
   m_cos[106]  =  13'b0011010101011;     //106pi/512
   m_sin[107]  =  13'b1101110001011;     //107pi/512
   m_cos[107]  =  13'b0011010100100;     //107pi/512
   m_sin[108]  =  13'b1101110000010;     //108pi/512
   m_cos[108]  =  13'b0011010011110;     //108pi/512
   m_sin[109]  =  13'b1101101111000;     //109pi/512
   m_cos[109]  =  13'b0011010011000;     //109pi/512
   m_sin[110]  =  13'b1101101101111;     //110pi/512
   m_cos[110]  =  13'b0011010010001;     //110pi/512
   m_sin[111]  =  13'b1101101100110;     //111pi/512
   m_cos[111]  =  13'b0011010001011;     //111pi/512
   m_sin[112]  =  13'b1101101011101;     //112pi/512
   m_cos[112]  =  13'b0011010000100;     //112pi/512
   m_sin[113]  =  13'b1101101010011;     //113pi/512
   m_cos[113]  =  13'b0011001111110;     //113pi/512
   m_sin[114]  =  13'b1101101001010;     //114pi/512
   m_cos[114]  =  13'b0011001110111;     //114pi/512
   m_sin[115]  =  13'b1101101000001;     //115pi/512
   m_cos[115]  =  13'b0011001110000;     //115pi/512
   m_sin[116]  =  13'b1101100111000;     //116pi/512
   m_cos[116]  =  13'b0011001101001;     //116pi/512
   m_sin[117]  =  13'b1101100101111;     //117pi/512
   m_cos[117]  =  13'b0011001100011;     //117pi/512
   m_sin[118]  =  13'b1101100100110;     //118pi/512
   m_cos[118]  =  13'b0011001011100;     //118pi/512
   m_sin[119]  =  13'b1101100011101;     //119pi/512
   m_cos[119]  =  13'b0011001010101;     //119pi/512
   m_sin[120]  =  13'b1101100010100;     //120pi/512
   m_cos[120]  =  13'b0011001001110;     //120pi/512
   m_sin[121]  =  13'b1101100001011;     //121pi/512
   m_cos[121]  =  13'b0011001000111;     //121pi/512
   m_sin[122]  =  13'b1101100000010;     //122pi/512
   m_cos[122]  =  13'b0011001000000;     //122pi/512
   m_sin[123]  =  13'b1101011111001;     //123pi/512
   m_cos[123]  =  13'b0011000111001;     //123pi/512
   m_sin[124]  =  13'b1101011110001;     //124pi/512
   m_cos[124]  =  13'b0011000110010;     //124pi/512
   m_sin[125]  =  13'b1101011101000;     //125pi/512
   m_cos[125]  =  13'b0011000101011;     //125pi/512
   m_sin[126]  =  13'b1101011011111;     //126pi/512
   m_cos[126]  =  13'b0011000100011;     //126pi/512
   m_sin[127]  =  13'b1101011010111;     //127pi/512
   m_cos[127]  =  13'b0011000011100;     //127pi/512
   m_sin[128]  =  13'b1101011001110;     //128pi/512
   m_cos[128]  =  13'b0011000010101;     //128pi/512
   m_sin[129]  =  13'b1101011000101;     //129pi/512
   m_cos[129]  =  13'b0011000001101;     //129pi/512
   m_sin[130]  =  13'b1101010111101;     //130pi/512
   m_cos[130]  =  13'b0011000000110;     //130pi/512
   m_sin[131]  =  13'b1101010110100;     //131pi/512
   m_cos[131]  =  13'b0010111111111;     //131pi/512
   m_sin[132]  =  13'b1101010101100;     //132pi/512
   m_cos[132]  =  13'b0010111110111;     //132pi/512
   m_sin[133]  =  13'b1101010100011;     //133pi/512
   m_cos[133]  =  13'b0010111101111;     //133pi/512
   m_sin[134]  =  13'b1101010011011;     //134pi/512
   m_cos[134]  =  13'b0010111101000;     //134pi/512
   m_sin[135]  =  13'b1101010010011;     //135pi/512
   m_cos[135]  =  13'b0010111100000;     //135pi/512
   m_sin[136]  =  13'b1101010001010;     //136pi/512
   m_cos[136]  =  13'b0010111011001;     //136pi/512
   m_sin[137]  =  13'b1101010000010;     //137pi/512
   m_cos[137]  =  13'b0010111010001;     //137pi/512
   m_sin[138]  =  13'b1101001111010;     //138pi/512
   m_cos[138]  =  13'b0010111001001;     //138pi/512
   m_sin[139]  =  13'b1101001110010;     //139pi/512
   m_cos[139]  =  13'b0010111000001;     //139pi/512
   m_sin[140]  =  13'b1101001101010;     //140pi/512
   m_cos[140]  =  13'b0010110111001;     //140pi/512
   m_sin[141]  =  13'b1101001100010;     //141pi/512
   m_cos[141]  =  13'b0010110110001;     //141pi/512
   m_sin[142]  =  13'b1101001011010;     //142pi/512
   m_cos[142]  =  13'b0010110101001;     //142pi/512
   m_sin[143]  =  13'b1101001010010;     //143pi/512
   m_cos[143]  =  13'b0010110100001;     //143pi/512
   m_sin[144]  =  13'b1101001001010;     //144pi/512
   m_cos[144]  =  13'b0010110011001;     //144pi/512
   m_sin[145]  =  13'b1101001000010;     //145pi/512
   m_cos[145]  =  13'b0010110010001;     //145pi/512
   m_sin[146]  =  13'b1101000111010;     //146pi/512
   m_cos[146]  =  13'b0010110001001;     //146pi/512
   m_sin[147]  =  13'b1101000110010;     //147pi/512
   m_cos[147]  =  13'b0010110000001;     //147pi/512
   m_sin[148]  =  13'b1101000101010;     //148pi/512
   m_cos[148]  =  13'b0010101111001;     //148pi/512
   m_sin[149]  =  13'b1101000100011;     //149pi/512
   m_cos[149]  =  13'b0010101110000;     //149pi/512
   m_sin[150]  =  13'b1101000011011;     //150pi/512
   m_cos[150]  =  13'b0010101101000;     //150pi/512
   m_sin[151]  =  13'b1101000010011;     //151pi/512
   m_cos[151]  =  13'b0010101100000;     //151pi/512
   m_sin[152]  =  13'b1101000001100;     //152pi/512
   m_cos[152]  =  13'b0010101010111;     //152pi/512
   m_sin[153]  =  13'b1101000000100;     //153pi/512
   m_cos[153]  =  13'b0010101001111;     //153pi/512
   m_sin[154]  =  13'b1100111111101;     //154pi/512
   m_cos[154]  =  13'b0010101000110;     //154pi/512
   m_sin[155]  =  13'b1100111110101;     //155pi/512
   m_cos[155]  =  13'b0010100111110;     //155pi/512
   m_sin[156]  =  13'b1100111101110;     //156pi/512
   m_cos[156]  =  13'b0010100110101;     //156pi/512
   m_sin[157]  =  13'b1100111100111;     //157pi/512
   m_cos[157]  =  13'b0010100101101;     //157pi/512
   m_sin[158]  =  13'b1100111011111;     //158pi/512
   m_cos[158]  =  13'b0010100100100;     //158pi/512
   m_sin[159]  =  13'b1100111011000;     //159pi/512
   m_cos[159]  =  13'b0010100011011;     //159pi/512
   m_sin[160]  =  13'b1100111010001;     //160pi/512
   m_cos[160]  =  13'b0010100010011;     //160pi/512
   m_sin[161]  =  13'b1100111001010;     //161pi/512
   m_cos[161]  =  13'b0010100001010;     //161pi/512
   m_sin[162]  =  13'b1100111000011;     //162pi/512
   m_cos[162]  =  13'b0010100000001;     //162pi/512
   m_sin[163]  =  13'b1100110111100;     //163pi/512
   m_cos[163]  =  13'b0010011111000;     //163pi/512
   m_sin[164]  =  13'b1100110110101;     //164pi/512
   m_cos[164]  =  13'b0010011101111;     //164pi/512
   m_sin[165]  =  13'b1100110101110;     //165pi/512
   m_cos[165]  =  13'b0010011100111;     //165pi/512
   m_sin[166]  =  13'b1100110100111;     //166pi/512
   m_cos[166]  =  13'b0010011011110;     //166pi/512
   m_sin[167]  =  13'b1100110100000;     //167pi/512
   m_cos[167]  =  13'b0010011010101;     //167pi/512
   m_sin[168]  =  13'b1100110011001;     //168pi/512
   m_cos[168]  =  13'b0010011001100;     //168pi/512
   m_sin[169]  =  13'b1100110010010;     //169pi/512
   m_cos[169]  =  13'b0010011000010;     //169pi/512
   m_sin[170]  =  13'b1100110001100;     //170pi/512
   m_cos[170]  =  13'b0010010111001;     //170pi/512
   m_sin[171]  =  13'b1100110000101;     //171pi/512
   m_cos[171]  =  13'b0010010110000;     //171pi/512
   m_sin[172]  =  13'b1100101111110;     //172pi/512
   m_cos[172]  =  13'b0010010100111;     //172pi/512
   m_sin[173]  =  13'b1100101111000;     //173pi/512
   m_cos[173]  =  13'b0010010011110;     //173pi/512
   m_sin[174]  =  13'b1100101110001;     //174pi/512
   m_cos[174]  =  13'b0010010010101;     //174pi/512
   m_sin[175]  =  13'b1100101101011;     //175pi/512
   m_cos[175]  =  13'b0010010001011;     //175pi/512
   m_sin[176]  =  13'b1100101100100;     //176pi/512
   m_cos[176]  =  13'b0010010000010;     //176pi/512
   m_sin[177]  =  13'b1100101011110;     //177pi/512
   m_cos[177]  =  13'b0010001111001;     //177pi/512
   m_sin[178]  =  13'b1100101011000;     //178pi/512
   m_cos[178]  =  13'b0010001101111;     //178pi/512
   m_sin[179]  =  13'b1100101010010;     //179pi/512
   m_cos[179]  =  13'b0010001100110;     //179pi/512
   m_sin[180]  =  13'b1100101001011;     //180pi/512
   m_cos[180]  =  13'b0010001011100;     //180pi/512
   m_sin[181]  =  13'b1100101000101;     //181pi/512
   m_cos[181]  =  13'b0010001010011;     //181pi/512
   m_sin[182]  =  13'b1100100111111;     //182pi/512
   m_cos[182]  =  13'b0010001001001;     //182pi/512
   m_sin[183]  =  13'b1100100111001;     //183pi/512
   m_cos[183]  =  13'b0010001000000;     //183pi/512
   m_sin[184]  =  13'b1100100110011;     //184pi/512
   m_cos[184]  =  13'b0010000110110;     //184pi/512
   m_sin[185]  =  13'b1100100101101;     //185pi/512
   m_cos[185]  =  13'b0010000101101;     //185pi/512
   m_sin[186]  =  13'b1100100100111;     //186pi/512
   m_cos[186]  =  13'b0010000100011;     //186pi/512
   m_sin[187]  =  13'b1100100100001;     //187pi/512
   m_cos[187]  =  13'b0010000011001;     //187pi/512
   m_sin[188]  =  13'b1100100011100;     //188pi/512
   m_cos[188]  =  13'b0010000001111;     //188pi/512
   m_sin[189]  =  13'b1100100010110;     //189pi/512
   m_cos[189]  =  13'b0010000000110;     //189pi/512
   m_sin[190]  =  13'b1100100010000;     //190pi/512
   m_cos[190]  =  13'b0001111111100;     //190pi/512
   m_sin[191]  =  13'b1100100001011;     //191pi/512
   m_cos[191]  =  13'b0001111110010;     //191pi/512
   m_sin[192]  =  13'b1100100000101;     //192pi/512
   m_cos[192]  =  13'b0001111101000;     //192pi/512
   m_sin[193]  =  13'b1100100000000;     //193pi/512
   m_cos[193]  =  13'b0001111011110;     //193pi/512
   m_sin[194]  =  13'b1100011111010;     //194pi/512
   m_cos[194]  =  13'b0001111010100;     //194pi/512
   m_sin[195]  =  13'b1100011110101;     //195pi/512
   m_cos[195]  =  13'b0001111001010;     //195pi/512
   m_sin[196]  =  13'b1100011101111;     //196pi/512
   m_cos[196]  =  13'b0001111000000;     //196pi/512
   m_sin[197]  =  13'b1100011101010;     //197pi/512
   m_cos[197]  =  13'b0001110110110;     //197pi/512
   m_sin[198]  =  13'b1100011100101;     //198pi/512
   m_cos[198]  =  13'b0001110101100;     //198pi/512
   m_sin[199]  =  13'b1100011100000;     //199pi/512
   m_cos[199]  =  13'b0001110100010;     //199pi/512
   m_sin[200]  =  13'b1100011011011;     //200pi/512
   m_cos[200]  =  13'b0001110011000;     //200pi/512
   m_sin[201]  =  13'b1100011010110;     //201pi/512
   m_cos[201]  =  13'b0001110001110;     //201pi/512
   m_sin[202]  =  13'b1100011010001;     //202pi/512
   m_cos[202]  =  13'b0001110000100;     //202pi/512
   m_sin[203]  =  13'b1100011001100;     //203pi/512
   m_cos[203]  =  13'b0001101111010;     //203pi/512
   m_sin[204]  =  13'b1100011000111;     //204pi/512
   m_cos[204]  =  13'b0001101110000;     //204pi/512
   m_sin[205]  =  13'b1100011000010;     //205pi/512
   m_cos[205]  =  13'b0001101100101;     //205pi/512
   m_sin[206]  =  13'b1100010111101;     //206pi/512
   m_cos[206]  =  13'b0001101011011;     //206pi/512
   m_sin[207]  =  13'b1100010111000;     //207pi/512
   m_cos[207]  =  13'b0001101010001;     //207pi/512
   m_sin[208]  =  13'b1100010110100;     //208pi/512
   m_cos[208]  =  13'b0001101000111;     //208pi/512
   m_sin[209]  =  13'b1100010101111;     //209pi/512
   m_cos[209]  =  13'b0001100111100;     //209pi/512
   m_sin[210]  =  13'b1100010101011;     //210pi/512
   m_cos[210]  =  13'b0001100110010;     //210pi/512
   m_sin[211]  =  13'b1100010100110;     //211pi/512
   m_cos[211]  =  13'b0001100101000;     //211pi/512
   m_sin[212]  =  13'b1100010100010;     //212pi/512
   m_cos[212]  =  13'b0001100011101;     //212pi/512
   m_sin[213]  =  13'b1100010011101;     //213pi/512
   m_cos[213]  =  13'b0001100010011;     //213pi/512
   m_sin[214]  =  13'b1100010011001;     //214pi/512
   m_cos[214]  =  13'b0001100001000;     //214pi/512
   m_sin[215]  =  13'b1100010010101;     //215pi/512
   m_cos[215]  =  13'b0001011111110;     //215pi/512
   m_sin[216]  =  13'b1100010010001;     //216pi/512
   m_cos[216]  =  13'b0001011110011;     //216pi/512
   m_sin[217]  =  13'b1100010001100;     //217pi/512
   m_cos[217]  =  13'b0001011101001;     //217pi/512
   m_sin[218]  =  13'b1100010001000;     //218pi/512
   m_cos[218]  =  13'b0001011011110;     //218pi/512
   m_sin[219]  =  13'b1100010000100;     //219pi/512
   m_cos[219]  =  13'b0001011010100;     //219pi/512
   m_sin[220]  =  13'b1100010000000;     //220pi/512
   m_cos[220]  =  13'b0001011001001;     //220pi/512
   m_sin[221]  =  13'b1100001111100;     //221pi/512
   m_cos[221]  =  13'b0001010111110;     //221pi/512
   m_sin[222]  =  13'b1100001111001;     //222pi/512
   m_cos[222]  =  13'b0001010110100;     //222pi/512
   m_sin[223]  =  13'b1100001110101;     //223pi/512
   m_cos[223]  =  13'b0001010101001;     //223pi/512
   m_sin[224]  =  13'b1100001110001;     //224pi/512
   m_cos[224]  =  13'b0001010011110;     //224pi/512
   m_sin[225]  =  13'b1100001101101;     //225pi/512
   m_cos[225]  =  13'b0001010010100;     //225pi/512
   m_sin[226]  =  13'b1100001101010;     //226pi/512
   m_cos[226]  =  13'b0001010001001;     //226pi/512
   m_sin[227]  =  13'b1100001100110;     //227pi/512
   m_cos[227]  =  13'b0001001111110;     //227pi/512
   m_sin[228]  =  13'b1100001100011;     //228pi/512
   m_cos[228]  =  13'b0001001110100;     //228pi/512
   m_sin[229]  =  13'b1100001011111;     //229pi/512
   m_cos[229]  =  13'b0001001101001;     //229pi/512
   m_sin[230]  =  13'b1100001011100;     //230pi/512
   m_cos[230]  =  13'b0001001011110;     //230pi/512
   m_sin[231]  =  13'b1100001011001;     //231pi/512
   m_cos[231]  =  13'b0001001010011;     //231pi/512
   m_sin[232]  =  13'b1100001010101;     //232pi/512
   m_cos[232]  =  13'b0001001001000;     //232pi/512
   m_sin[233]  =  13'b1100001010010;     //233pi/512
   m_cos[233]  =  13'b0001000111110;     //233pi/512
   m_sin[234]  =  13'b1100001001111;     //234pi/512
   m_cos[234]  =  13'b0001000110011;     //234pi/512
   m_sin[235]  =  13'b1100001001100;     //235pi/512
   m_cos[235]  =  13'b0001000101000;     //235pi/512
   m_sin[236]  =  13'b1100001001001;     //236pi/512
   m_cos[236]  =  13'b0001000011101;     //236pi/512
   m_sin[237]  =  13'b1100001000110;     //237pi/512
   m_cos[237]  =  13'b0001000010010;     //237pi/512
   m_sin[238]  =  13'b1100001000011;     //238pi/512
   m_cos[238]  =  13'b0001000000111;     //238pi/512
   m_sin[239]  =  13'b1100001000000;     //239pi/512
   m_cos[239]  =  13'b0000111111100;     //239pi/512
   m_sin[240]  =  13'b1100000111101;     //240pi/512
   m_cos[240]  =  13'b0000111110001;     //240pi/512
   m_sin[241]  =  13'b1100000111011;     //241pi/512
   m_cos[241]  =  13'b0000111100110;     //241pi/512
   m_sin[242]  =  13'b1100000111000;     //242pi/512
   m_cos[242]  =  13'b0000111011011;     //242pi/512
   m_sin[243]  =  13'b1100000110101;     //243pi/512
   m_cos[243]  =  13'b0000111010000;     //243pi/512
   m_sin[244]  =  13'b1100000110011;     //244pi/512
   m_cos[244]  =  13'b0000111000101;     //244pi/512
   m_sin[245]  =  13'b1100000110000;     //245pi/512
   m_cos[245]  =  13'b0000110111010;     //245pi/512
   m_sin[246]  =  13'b1100000101110;     //246pi/512
   m_cos[246]  =  13'b0000110101111;     //246pi/512
   m_sin[247]  =  13'b1100000101100;     //247pi/512
   m_cos[247]  =  13'b0000110100100;     //247pi/512
   m_sin[248]  =  13'b1100000101001;     //248pi/512
   m_cos[248]  =  13'b0000110011001;     //248pi/512
   m_sin[249]  =  13'b1100000100111;     //249pi/512
   m_cos[249]  =  13'b0000110001110;     //249pi/512
   m_sin[250]  =  13'b1100000100101;     //250pi/512
   m_cos[250]  =  13'b0000110000011;     //250pi/512
   m_sin[251]  =  13'b1100000100011;     //251pi/512
   m_cos[251]  =  13'b0000101111000;     //251pi/512
   m_sin[252]  =  13'b1100000100001;     //252pi/512
   m_cos[252]  =  13'b0000101101100;     //252pi/512
   m_sin[253]  =  13'b1100000011111;     //253pi/512
   m_cos[253]  =  13'b0000101100001;     //253pi/512
   m_sin[254]  =  13'b1100000011101;     //254pi/512
   m_cos[254]  =  13'b0000101010110;     //254pi/512
   m_sin[255]  =  13'b1100000011011;     //255pi/512
   m_cos[255]  =  13'b0000101001011;     //255pi/512
   m_sin[256]  =  13'b1100000011001;     //256pi/512
   m_cos[256]  =  13'b0000101000000;     //256pi/512
   m_sin[257]  =  13'b1100000010111;     //257pi/512
   m_cos[257]  =  13'b0000100110101;     //257pi/512
   m_sin[258]  =  13'b1100000010110;     //258pi/512
   m_cos[258]  =  13'b0000100101010;     //258pi/512
   m_sin[259]  =  13'b1100000010100;     //259pi/512
   m_cos[259]  =  13'b0000100011110;     //259pi/512
   m_sin[260]  =  13'b1100000010011;     //260pi/512
   m_cos[260]  =  13'b0000100010011;     //260pi/512
   m_sin[261]  =  13'b1100000010001;     //261pi/512
   m_cos[261]  =  13'b0000100001000;     //261pi/512
   m_sin[262]  =  13'b1100000010000;     //262pi/512
   m_cos[262]  =  13'b0000011111101;     //262pi/512
   m_sin[263]  =  13'b1100000001110;     //263pi/512
   m_cos[263]  =  13'b0000011110001;     //263pi/512
   m_sin[264]  =  13'b1100000001101;     //264pi/512
   m_cos[264]  =  13'b0000011100110;     //264pi/512
   m_sin[265]  =  13'b1100000001100;     //265pi/512
   m_cos[265]  =  13'b0000011011011;     //265pi/512
   m_sin[266]  =  13'b1100000001011;     //266pi/512
   m_cos[266]  =  13'b0000011010000;     //266pi/512
   m_sin[267]  =  13'b1100000001001;     //267pi/512
   m_cos[267]  =  13'b0000011000100;     //267pi/512
   m_sin[268]  =  13'b1100000001000;     //268pi/512
   m_cos[268]  =  13'b0000010111001;     //268pi/512
   m_sin[269]  =  13'b1100000000111;     //269pi/512
   m_cos[269]  =  13'b0000010101110;     //269pi/512
   m_sin[270]  =  13'b1100000000111;     //270pi/512
   m_cos[270]  =  13'b0000010100011;     //270pi/512
   m_sin[271]  =  13'b1100000000110;     //271pi/512
   m_cos[271]  =  13'b0000010010111;     //271pi/512
   m_sin[272]  =  13'b1100000000101;     //272pi/512
   m_cos[272]  =  13'b0000010001100;     //272pi/512
   m_sin[273]  =  13'b1100000000100;     //273pi/512
   m_cos[273]  =  13'b0000010000001;     //273pi/512
   m_sin[274]  =  13'b1100000000011;     //274pi/512
   m_cos[274]  =  13'b0000001110110;     //274pi/512
   m_sin[275]  =  13'b1100000000011;     //275pi/512
   m_cos[275]  =  13'b0000001101010;     //275pi/512
   m_sin[276]  =  13'b1100000000010;     //276pi/512
   m_cos[276]  =  13'b0000001011111;     //276pi/512
   m_sin[277]  =  13'b1100000000010;     //277pi/512
   m_cos[277]  =  13'b0000001010100;     //277pi/512
   m_sin[278]  =  13'b1100000000001;     //278pi/512
   m_cos[278]  =  13'b0000001001000;     //278pi/512
   m_sin[279]  =  13'b1100000000001;     //279pi/512
   m_cos[279]  =  13'b0000000111101;     //279pi/512
   m_sin[280]  =  13'b1100000000001;     //280pi/512
   m_cos[280]  =  13'b0000000110010;     //280pi/512
   m_sin[281]  =  13'b1100000000000;     //281pi/512
   m_cos[281]  =  13'b0000000100110;     //281pi/512
   m_sin[282]  =  13'b1100000000000;     //282pi/512
   m_cos[282]  =  13'b0000000011011;     //282pi/512
   m_sin[283]  =  13'b1100000000000;     //283pi/512
   m_cos[283]  =  13'b0000000010000;     //283pi/512
   m_sin[284]  =  13'b1100000000000;     //284pi/512
   m_cos[284]  =  13'b0000000000101;     //284pi/512
   m_sin[285]  =  13'b1100000000000;     //285pi/512
   m_cos[285]  =  13'b1111111111010;     //285pi/512
   m_sin[286]  =  13'b1100000000000;     //286pi/512
   m_cos[286]  =  13'b1111111101110;     //286pi/512
   m_sin[287]  =  13'b1100000000000;     //287pi/512
   m_cos[287]  =  13'b1111111100011;     //287pi/512
   m_sin[288]  =  13'b1100000000000;     //288pi/512
   m_cos[288]  =  13'b1111111011000;     //288pi/512
   m_sin[289]  =  13'b1100000000001;     //289pi/512
   m_cos[289]  =  13'b1111111001100;     //289pi/512
   m_sin[290]  =  13'b1100000000001;     //290pi/512
   m_cos[290]  =  13'b1111111000001;     //290pi/512
   m_sin[291]  =  13'b1100000000001;     //291pi/512
   m_cos[291]  =  13'b1111110110110;     //291pi/512
   m_sin[292]  =  13'b1100000000010;     //292pi/512
   m_cos[292]  =  13'b1111110101011;     //292pi/512
   m_sin[293]  =  13'b1100000000010;     //293pi/512
   m_cos[293]  =  13'b1111110011111;     //293pi/512
   m_sin[294]  =  13'b1100000000011;     //294pi/512
   m_cos[294]  =  13'b1111110010100;     //294pi/512
   m_sin[295]  =  13'b1100000000011;     //295pi/512
   m_cos[295]  =  13'b1111110001001;     //295pi/512
   m_sin[296]  =  13'b1100000000100;     //296pi/512
   m_cos[296]  =  13'b1111101111101;     //296pi/512
   m_sin[297]  =  13'b1100000000101;     //297pi/512
   m_cos[297]  =  13'b1111101110010;     //297pi/512
   m_sin[298]  =  13'b1100000000110;     //298pi/512
   m_cos[298]  =  13'b1111101100111;     //298pi/512
   m_sin[299]  =  13'b1100000000111;     //299pi/512
   m_cos[299]  =  13'b1111101011100;     //299pi/512
   m_sin[300]  =  13'b1100000001000;     //300pi/512
   m_cos[300]  =  13'b1111101010000;     //300pi/512
   m_sin[301]  =  13'b1100000001001;     //301pi/512
   m_cos[301]  =  13'b1111101000101;     //301pi/512
   m_sin[302]  =  13'b1100000001010;     //302pi/512
   m_cos[302]  =  13'b1111100111010;     //302pi/512
   m_sin[303]  =  13'b1100000001011;     //303pi/512
   m_cos[303]  =  13'b1111100101111;     //303pi/512
   m_sin[304]  =  13'b1100000001100;     //304pi/512
   m_cos[304]  =  13'b1111100100011;     //304pi/512
   m_sin[305]  =  13'b1100000001101;     //305pi/512
   m_cos[305]  =  13'b1111100011000;     //305pi/512
   m_sin[306]  =  13'b1100000001110;     //306pi/512
   m_cos[306]  =  13'b1111100001101;     //306pi/512
   m_sin[307]  =  13'b1100000010000;     //307pi/512
   m_cos[307]  =  13'b1111100000010;     //307pi/512
   m_sin[308]  =  13'b1100000010001;     //308pi/512
   m_cos[308]  =  13'b1111011110110;     //308pi/512
   m_sin[309]  =  13'b1100000010011;     //309pi/512
   m_cos[309]  =  13'b1111011101011;     //309pi/512
   m_sin[310]  =  13'b1100000010100;     //310pi/512
   m_cos[310]  =  13'b1111011100000;     //310pi/512
   m_sin[311]  =  13'b1100000010110;     //311pi/512
   m_cos[311]  =  13'b1111011010101;     //311pi/512
   m_sin[312]  =  13'b1100000011000;     //312pi/512
   m_cos[312]  =  13'b1111011001010;     //312pi/512
   m_sin[313]  =  13'b1100000011001;     //313pi/512
   m_cos[313]  =  13'b1111010111110;     //313pi/512
   m_sin[314]  =  13'b1100000011011;     //314pi/512
   m_cos[314]  =  13'b1111010110011;     //314pi/512
   m_sin[315]  =  13'b1100000011101;     //315pi/512
   m_cos[315]  =  13'b1111010101000;     //315pi/512
   m_sin[316]  =  13'b1100000011111;     //316pi/512
   m_cos[316]  =  13'b1111010011101;     //316pi/512
   m_sin[317]  =  13'b1100000100001;     //317pi/512
   m_cos[317]  =  13'b1111010010010;     //317pi/512
   m_sin[318]  =  13'b1100000100011;     //318pi/512
   m_cos[318]  =  13'b1111010000111;     //318pi/512
   m_sin[319]  =  13'b1100000100101;     //319pi/512
   m_cos[319]  =  13'b1111001111100;     //319pi/512
   m_sin[320]  =  13'b1100000100111;     //320pi/512
   m_cos[320]  =  13'b1111001110000;     //320pi/512
   m_sin[321]  =  13'b1100000101010;     //321pi/512
   m_cos[321]  =  13'b1111001100101;     //321pi/512
   m_sin[322]  =  13'b1100000101100;     //322pi/512
   m_cos[322]  =  13'b1111001011010;     //322pi/512
   m_sin[323]  =  13'b1100000101110;     //323pi/512
   m_cos[323]  =  13'b1111001001111;     //323pi/512
   m_sin[324]  =  13'b1100000110001;     //324pi/512
   m_cos[324]  =  13'b1111001000100;     //324pi/512
   m_sin[325]  =  13'b1100000110011;     //325pi/512
   m_cos[325]  =  13'b1111000111001;     //325pi/512
   m_sin[326]  =  13'b1100000110110;     //326pi/512
   m_cos[326]  =  13'b1111000101110;     //326pi/512
   m_sin[327]  =  13'b1100000111000;     //327pi/512
   m_cos[327]  =  13'b1111000100011;     //327pi/512
   m_sin[328]  =  13'b1100000111011;     //328pi/512
   m_cos[328]  =  13'b1111000011000;     //328pi/512
   m_sin[329]  =  13'b1100000111110;     //329pi/512
   m_cos[329]  =  13'b1111000001101;     //329pi/512
   m_sin[330]  =  13'b1100001000000;     //330pi/512
   m_cos[330]  =  13'b1111000000010;     //330pi/512
   m_sin[331]  =  13'b1100001000011;     //331pi/512
   m_cos[331]  =  13'b1110111110111;     //331pi/512
   m_sin[332]  =  13'b1100001000110;     //332pi/512
   m_cos[332]  =  13'b1110111101100;     //332pi/512
   m_sin[333]  =  13'b1100001001001;     //333pi/512
   m_cos[333]  =  13'b1110111100001;     //333pi/512
   m_sin[334]  =  13'b1100001001100;     //334pi/512
   m_cos[334]  =  13'b1110111010111;     //334pi/512
   m_sin[335]  =  13'b1100001001111;     //335pi/512
   m_cos[335]  =  13'b1110111001100;     //335pi/512
   m_sin[336]  =  13'b1100001010010;     //336pi/512
   m_cos[336]  =  13'b1110111000001;     //336pi/512
   m_sin[337]  =  13'b1100001010110;     //337pi/512
   m_cos[337]  =  13'b1110110110110;     //337pi/512
   m_sin[338]  =  13'b1100001011001;     //338pi/512
   m_cos[338]  =  13'b1110110101011;     //338pi/512
   m_sin[339]  =  13'b1100001011100;     //339pi/512
   m_cos[339]  =  13'b1110110100000;     //339pi/512
   m_sin[340]  =  13'b1100001100000;     //340pi/512
   m_cos[340]  =  13'b1110110010101;     //340pi/512
   m_sin[341]  =  13'b1100001100011;     //341pi/512
   m_cos[341]  =  13'b1110110001011;     //341pi/512
   m_sin[342]  =  13'b1100001100111;     //342pi/512
   m_cos[342]  =  13'b1110110000000;     //342pi/512
   m_sin[343]  =  13'b1100001101010;     //343pi/512
   m_cos[343]  =  13'b1110101110101;     //343pi/512
   m_sin[344]  =  13'b1100001101110;     //344pi/512
   m_cos[344]  =  13'b1110101101011;     //344pi/512
   m_sin[345]  =  13'b1100001110001;     //345pi/512
   m_cos[345]  =  13'b1110101100000;     //345pi/512
   m_sin[346]  =  13'b1100001110101;     //346pi/512
   m_cos[346]  =  13'b1110101010101;     //346pi/512
   m_sin[347]  =  13'b1100001111001;     //347pi/512
   m_cos[347]  =  13'b1110101001011;     //347pi/512
   m_sin[348]  =  13'b1100001111101;     //348pi/512
   m_cos[348]  =  13'b1110101000000;     //348pi/512
   m_sin[349]  =  13'b1100010000001;     //349pi/512
   m_cos[349]  =  13'b1110100110101;     //349pi/512
   m_sin[350]  =  13'b1100010000101;     //350pi/512
   m_cos[350]  =  13'b1110100101011;     //350pi/512
   m_sin[351]  =  13'b1100010001001;     //351pi/512
   m_cos[351]  =  13'b1110100100000;     //351pi/512
   m_sin[352]  =  13'b1100010001101;     //352pi/512
   m_cos[352]  =  13'b1110100010110;     //352pi/512
   m_sin[353]  =  13'b1100010010001;     //353pi/512
   m_cos[353]  =  13'b1110100001011;     //353pi/512
   m_sin[354]  =  13'b1100010010101;     //354pi/512
   m_cos[354]  =  13'b1110100000001;     //354pi/512
   m_sin[355]  =  13'b1100010011001;     //355pi/512
   m_cos[355]  =  13'b1110011110110;     //355pi/512
   m_sin[356]  =  13'b1100010011110;     //356pi/512
   m_cos[356]  =  13'b1110011101100;     //356pi/512
   m_sin[357]  =  13'b1100010100010;     //357pi/512
   m_cos[357]  =  13'b1110011100001;     //357pi/512
   m_sin[358]  =  13'b1100010100111;     //358pi/512
   m_cos[358]  =  13'b1110011010111;     //358pi/512
   m_sin[359]  =  13'b1100010101011;     //359pi/512
   m_cos[359]  =  13'b1110011001100;     //359pi/512
   m_sin[360]  =  13'b1100010110000;     //360pi/512
   m_cos[360]  =  13'b1110011000010;     //360pi/512
   m_sin[361]  =  13'b1100010110100;     //361pi/512
   m_cos[361]  =  13'b1110010111000;     //361pi/512
   m_sin[362]  =  13'b1100010111001;     //362pi/512
   m_cos[362]  =  13'b1110010101101;     //362pi/512
   m_sin[363]  =  13'b1100010111110;     //363pi/512
   m_cos[363]  =  13'b1110010100011;     //363pi/512
   m_sin[364]  =  13'b1100011000010;     //364pi/512
   m_cos[364]  =  13'b1110010011001;     //364pi/512
   m_sin[365]  =  13'b1100011000111;     //365pi/512
   m_cos[365]  =  13'b1110010001111;     //365pi/512
   m_sin[366]  =  13'b1100011001100;     //366pi/512
   m_cos[366]  =  13'b1110010000100;     //366pi/512
   m_sin[367]  =  13'b1100011010001;     //367pi/512
   m_cos[367]  =  13'b1110001111010;     //367pi/512
   m_sin[368]  =  13'b1100011010110;     //368pi/512
   m_cos[368]  =  13'b1110001110000;     //368pi/512
   m_sin[369]  =  13'b1100011011011;     //369pi/512
   m_cos[369]  =  13'b1110001100110;     //369pi/512
   m_sin[370]  =  13'b1100011100000;     //370pi/512
   m_cos[370]  =  13'b1110001011100;     //370pi/512
   m_sin[371]  =  13'b1100011100110;     //371pi/512
   m_cos[371]  =  13'b1110001010010;     //371pi/512
   m_sin[372]  =  13'b1100011101011;     //372pi/512
   m_cos[372]  =  13'b1110001001000;     //372pi/512
   m_sin[373]  =  13'b1100011110000;     //373pi/512
   m_cos[373]  =  13'b1110000111110;     //373pi/512
   m_sin[374]  =  13'b1100011110101;     //374pi/512
   m_cos[374]  =  13'b1110000110100;     //374pi/512
   m_sin[375]  =  13'b1100011111011;     //375pi/512
   m_cos[375]  =  13'b1110000101010;     //375pi/512
   m_sin[376]  =  13'b1100100000000;     //376pi/512
   m_cos[376]  =  13'b1110000100000;     //376pi/512
   m_sin[377]  =  13'b1100100000110;     //377pi/512
   m_cos[377]  =  13'b1110000010110;     //377pi/512
   m_sin[378]  =  13'b1100100001011;     //378pi/512
   m_cos[378]  =  13'b1110000001100;     //378pi/512
   m_sin[379]  =  13'b1100100010001;     //379pi/512
   m_cos[379]  =  13'b1110000000011;     //379pi/512
   m_sin[380]  =  13'b1100100010111;     //380pi/512
   m_cos[380]  =  13'b1101111111001;     //380pi/512
   m_sin[381]  =  13'b1100100011100;     //381pi/512
   m_cos[381]  =  13'b1101111101111;     //381pi/512
   m_sin[382]  =  13'b1100100100010;     //382pi/512
   m_cos[382]  =  13'b1101111100101;     //382pi/512
   m_sin[383]  =  13'b1100100101000;     //383pi/512
   m_cos[383]  =  13'b1101111011100;     //383pi/512
   m_sin[384]  =  13'b1100100101110;     //384pi/512
   m_cos[384]  =  13'b1101111010010;     //384pi/512
   m_sin[385]  =  13'b1100100110100;     //385pi/512
   m_cos[385]  =  13'b1101111001000;     //385pi/512
   m_sin[386]  =  13'b1100100111010;     //386pi/512
   m_cos[386]  =  13'b1101110111111;     //386pi/512
   m_sin[387]  =  13'b1100101000000;     //387pi/512
   m_cos[387]  =  13'b1101110110101;     //387pi/512
   m_sin[388]  =  13'b1100101000110;     //388pi/512
   m_cos[388]  =  13'b1101110101100;     //388pi/512
   m_sin[389]  =  13'b1100101001100;     //389pi/512
   m_cos[389]  =  13'b1101110100010;     //389pi/512
   m_sin[390]  =  13'b1100101010010;     //390pi/512
   m_cos[390]  =  13'b1101110011001;     //390pi/512
   m_sin[391]  =  13'b1100101011000;     //391pi/512
   m_cos[391]  =  13'b1101110001111;     //391pi/512
   m_sin[392]  =  13'b1100101011111;     //392pi/512
   m_cos[392]  =  13'b1101110000110;     //392pi/512
   m_sin[393]  =  13'b1100101100101;     //393pi/512
   m_cos[393]  =  13'b1101101111100;     //393pi/512
   m_sin[394]  =  13'b1100101101100;     //394pi/512
   m_cos[394]  =  13'b1101101110011;     //394pi/512
   m_sin[395]  =  13'b1100101110010;     //395pi/512
   m_cos[395]  =  13'b1101101101010;     //395pi/512
   m_sin[396]  =  13'b1100101111000;     //396pi/512
   m_cos[396]  =  13'b1101101100001;     //396pi/512
   m_sin[397]  =  13'b1100101111111;     //397pi/512
   m_cos[397]  =  13'b1101101010111;     //397pi/512
   m_sin[398]  =  13'b1100110000110;     //398pi/512
   m_cos[398]  =  13'b1101101001110;     //398pi/512
   m_sin[399]  =  13'b1100110001100;     //399pi/512
   m_cos[399]  =  13'b1101101000101;     //399pi/512
   m_sin[400]  =  13'b1100110010011;     //400pi/512
   m_cos[400]  =  13'b1101100111100;     //400pi/512
   m_sin[401]  =  13'b1100110011010;     //401pi/512
   m_cos[401]  =  13'b1101100110011;     //401pi/512
   m_sin[402]  =  13'b1100110100001;     //402pi/512
   m_cos[402]  =  13'b1101100101010;     //402pi/512
   m_sin[403]  =  13'b1100110100111;     //403pi/512
   m_cos[403]  =  13'b1101100100001;     //403pi/512
   m_sin[404]  =  13'b1100110101110;     //404pi/512
   m_cos[404]  =  13'b1101100011000;     //404pi/512
   m_sin[405]  =  13'b1100110110101;     //405pi/512
   m_cos[405]  =  13'b1101100001111;     //405pi/512
   m_sin[406]  =  13'b1100110111100;     //406pi/512
   m_cos[406]  =  13'b1101100000110;     //406pi/512
   m_sin[407]  =  13'b1100111000011;     //407pi/512
   m_cos[407]  =  13'b1101011111101;     //407pi/512
   m_sin[408]  =  13'b1100111001011;     //408pi/512
   m_cos[408]  =  13'b1101011110101;     //408pi/512
   m_sin[409]  =  13'b1100111010010;     //409pi/512
   m_cos[409]  =  13'b1101011101100;     //409pi/512
   m_sin[410]  =  13'b1100111011001;     //410pi/512
   m_cos[410]  =  13'b1101011100011;     //410pi/512
   m_sin[411]  =  13'b1100111100000;     //411pi/512
   m_cos[411]  =  13'b1101011011010;     //411pi/512
   m_sin[412]  =  13'b1100111100111;     //412pi/512
   m_cos[412]  =  13'b1101011010010;     //412pi/512
   m_sin[413]  =  13'b1100111101111;     //413pi/512
   m_cos[413]  =  13'b1101011001001;     //413pi/512
   m_sin[414]  =  13'b1100111110110;     //414pi/512
   m_cos[414]  =  13'b1101011000001;     //414pi/512
   m_sin[415]  =  13'b1100111111110;     //415pi/512
   m_cos[415]  =  13'b1101010111000;     //415pi/512
   m_sin[416]  =  13'b1101000000101;     //416pi/512
   m_cos[416]  =  13'b1101010110000;     //416pi/512
   m_sin[417]  =  13'b1101000001101;     //417pi/512
   m_cos[417]  =  13'b1101010100111;     //417pi/512
   m_sin[418]  =  13'b1101000010100;     //418pi/512
   m_cos[418]  =  13'b1101010011111;     //418pi/512
   m_sin[419]  =  13'b1101000011100;     //419pi/512
   m_cos[419]  =  13'b1101010010110;     //419pi/512
   m_sin[420]  =  13'b1101000100100;     //420pi/512
   m_cos[420]  =  13'b1101010001110;     //420pi/512
   m_sin[421]  =  13'b1101000101011;     //421pi/512
   m_cos[421]  =  13'b1101010000110;     //421pi/512
   m_sin[422]  =  13'b1101000110011;     //422pi/512
   m_cos[422]  =  13'b1101001111110;     //422pi/512
   m_sin[423]  =  13'b1101000111011;     //423pi/512
   m_cos[423]  =  13'b1101001110101;     //423pi/512
   m_sin[424]  =  13'b1101001000011;     //424pi/512
   m_cos[424]  =  13'b1101001101101;     //424pi/512
   m_sin[425]  =  13'b1101001001011;     //425pi/512
   m_cos[425]  =  13'b1101001100101;     //425pi/512
   m_sin[426]  =  13'b1101001010011;     //426pi/512
   m_cos[426]  =  13'b1101001011101;     //426pi/512
   m_sin[427]  =  13'b1101001011011;     //427pi/512
   m_cos[427]  =  13'b1101001010101;     //427pi/512
   m_sin[428]  =  13'b1101001100011;     //428pi/512
   m_cos[428]  =  13'b1101001001101;     //428pi/512
   m_sin[429]  =  13'b1101001101011;     //429pi/512
   m_cos[429]  =  13'b1101001000101;     //429pi/512
   m_sin[430]  =  13'b1101001110011;     //430pi/512
   m_cos[430]  =  13'b1101000111101;     //430pi/512
   m_sin[431]  =  13'b1101001111011;     //431pi/512
   m_cos[431]  =  13'b1101000110110;     //431pi/512
   m_sin[432]  =  13'b1101010000011;     //432pi/512
   m_cos[432]  =  13'b1101000101110;     //432pi/512
   m_sin[433]  =  13'b1101010001011;     //433pi/512
   m_cos[433]  =  13'b1101000100110;     //433pi/512
   m_sin[434]  =  13'b1101010010100;     //434pi/512
   m_cos[434]  =  13'b1101000011110;     //434pi/512
   m_sin[435]  =  13'b1101010011100;     //435pi/512
   m_cos[435]  =  13'b1101000010111;     //435pi/512
   m_sin[436]  =  13'b1101010100100;     //436pi/512
   m_cos[436]  =  13'b1101000001111;     //436pi/512
   m_sin[437]  =  13'b1101010101101;     //437pi/512
   m_cos[437]  =  13'b1101000001000;     //437pi/512
   m_sin[438]  =  13'b1101010110101;     //438pi/512
   m_cos[438]  =  13'b1101000000000;     //438pi/512
   m_sin[439]  =  13'b1101010111110;     //439pi/512
   m_cos[439]  =  13'b1100111111001;     //439pi/512
   m_sin[440]  =  13'b1101011000110;     //440pi/512
   m_cos[440]  =  13'b1100111110001;     //440pi/512
   m_sin[441]  =  13'b1101011001111;     //441pi/512
   m_cos[441]  =  13'b1100111101010;     //441pi/512
   m_sin[442]  =  13'b1101011011000;     //442pi/512
   m_cos[442]  =  13'b1100111100011;     //442pi/512
   m_sin[443]  =  13'b1101011100000;     //443pi/512
   m_cos[443]  =  13'b1100111011011;     //443pi/512
   m_sin[444]  =  13'b1101011101001;     //444pi/512
   m_cos[444]  =  13'b1100111010100;     //444pi/512
   m_sin[445]  =  13'b1101011110010;     //445pi/512
   m_cos[445]  =  13'b1100111001101;     //445pi/512
   m_sin[446]  =  13'b1101011111010;     //446pi/512
   m_cos[446]  =  13'b1100111000110;     //446pi/512
   m_sin[447]  =  13'b1101100000011;     //447pi/512
   m_cos[447]  =  13'b1100110111111;     //447pi/512
   m_sin[448]  =  13'b1101100001100;     //448pi/512
   m_cos[448]  =  13'b1100110111000;     //448pi/512
   m_sin[449]  =  13'b1101100010101;     //449pi/512
   m_cos[449]  =  13'b1100110110001;     //449pi/512
   m_sin[450]  =  13'b1101100011110;     //450pi/512
   m_cos[450]  =  13'b1100110101010;     //450pi/512
   m_sin[451]  =  13'b1101100100111;     //451pi/512
   m_cos[451]  =  13'b1100110100011;     //451pi/512
   m_sin[452]  =  13'b1101100110000;     //452pi/512
   m_cos[452]  =  13'b1100110011100;     //452pi/512
   m_sin[453]  =  13'b1101100111001;     //453pi/512
   m_cos[453]  =  13'b1100110010101;     //453pi/512
   m_sin[454]  =  13'b1101101000010;     //454pi/512
   m_cos[454]  =  13'b1100110001111;     //454pi/512
   m_sin[455]  =  13'b1101101001011;     //455pi/512
   m_cos[455]  =  13'b1100110001000;     //455pi/512
   m_sin[456]  =  13'b1101101010100;     //456pi/512
   m_cos[456]  =  13'b1100110000001;     //456pi/512
   m_sin[457]  =  13'b1101101011110;     //457pi/512
   m_cos[457]  =  13'b1100101111011;     //457pi/512
   m_sin[458]  =  13'b1101101100111;     //458pi/512
   m_cos[458]  =  13'b1100101110100;     //458pi/512
   m_sin[459]  =  13'b1101101110000;     //459pi/512
   m_cos[459]  =  13'b1100101101110;     //459pi/512
   m_sin[460]  =  13'b1101101111001;     //460pi/512
   m_cos[460]  =  13'b1100101100111;     //460pi/512
   m_sin[461]  =  13'b1101110000011;     //461pi/512
   m_cos[461]  =  13'b1100101100001;     //461pi/512
   m_sin[462]  =  13'b1101110001100;     //462pi/512
   m_cos[462]  =  13'b1100101011011;     //462pi/512
   m_sin[463]  =  13'b1101110010110;     //463pi/512
   m_cos[463]  =  13'b1100101010100;     //463pi/512
   m_sin[464]  =  13'b1101110011111;     //464pi/512
   m_cos[464]  =  13'b1100101001110;     //464pi/512
   m_sin[465]  =  13'b1101110101000;     //465pi/512
   m_cos[465]  =  13'b1100101001000;     //465pi/512
   m_sin[466]  =  13'b1101110110010;     //466pi/512
   m_cos[466]  =  13'b1100101000010;     //466pi/512
   m_sin[467]  =  13'b1101110111100;     //467pi/512
   m_cos[467]  =  13'b1100100111100;     //467pi/512
   m_sin[468]  =  13'b1101111000101;     //468pi/512
   m_cos[468]  =  13'b1100100110110;     //468pi/512
   m_sin[469]  =  13'b1101111001111;     //469pi/512
   m_cos[469]  =  13'b1100100110000;     //469pi/512
   m_sin[470]  =  13'b1101111011000;     //470pi/512
   m_cos[470]  =  13'b1100100101010;     //470pi/512
   m_sin[471]  =  13'b1101111100010;     //471pi/512
   m_cos[471]  =  13'b1100100100100;     //471pi/512
   m_sin[472]  =  13'b1101111101100;     //472pi/512
   m_cos[472]  =  13'b1100100011110;     //472pi/512
   m_sin[473]  =  13'b1101111110101;     //473pi/512
   m_cos[473]  =  13'b1100100011000;     //473pi/512
   m_sin[474]  =  13'b1101111111111;     //474pi/512
   m_cos[474]  =  13'b1100100010011;     //474pi/512
   m_sin[475]  =  13'b1110000001001;     //475pi/512
   m_cos[475]  =  13'b1100100001101;     //475pi/512
   m_sin[476]  =  13'b1110000010011;     //476pi/512
   m_cos[476]  =  13'b1100100001000;     //476pi/512
   m_sin[477]  =  13'b1110000011101;     //477pi/512
   m_cos[477]  =  13'b1100100000010;     //477pi/512
   m_sin[478]  =  13'b1110000100111;     //478pi/512
   m_cos[478]  =  13'b1100011111101;     //478pi/512
   m_sin[479]  =  13'b1110000110001;     //479pi/512
   m_cos[479]  =  13'b1100011110111;     //479pi/512
   m_sin[480]  =  13'b1110000111011;     //480pi/512
   m_cos[480]  =  13'b1100011110010;     //480pi/512
   m_sin[481]  =  13'b1110001000101;     //481pi/512
   m_cos[481]  =  13'b1100011101101;     //481pi/512
   m_sin[482]  =  13'b1110001001111;     //482pi/512
   m_cos[482]  =  13'b1100011100111;     //482pi/512
   m_sin[483]  =  13'b1110001011001;     //483pi/512
   m_cos[483]  =  13'b1100011100010;     //483pi/512
   m_sin[484]  =  13'b1110001100011;     //484pi/512
   m_cos[484]  =  13'b1100011011101;     //484pi/512
   m_sin[485]  =  13'b1110001101101;     //485pi/512
   m_cos[485]  =  13'b1100011011000;     //485pi/512
   m_sin[486]  =  13'b1110001110111;     //486pi/512
   m_cos[486]  =  13'b1100011010011;     //486pi/512
   m_sin[487]  =  13'b1110010000001;     //487pi/512
   m_cos[487]  =  13'b1100011001110;     //487pi/512
   m_sin[488]  =  13'b1110010001011;     //488pi/512
   m_cos[488]  =  13'b1100011001001;     //488pi/512
   m_sin[489]  =  13'b1110010010110;     //489pi/512
   m_cos[489]  =  13'b1100011000100;     //489pi/512
   m_sin[490]  =  13'b1110010100000;     //490pi/512
   m_cos[490]  =  13'b1100010111111;     //490pi/512
   m_sin[491]  =  13'b1110010101010;     //491pi/512
   m_cos[491]  =  13'b1100010111011;     //491pi/512
   m_sin[492]  =  13'b1110010110100;     //492pi/512
   m_cos[492]  =  13'b1100010110110;     //492pi/512
   m_sin[493]  =  13'b1110010111111;     //493pi/512
   m_cos[493]  =  13'b1100010110001;     //493pi/512
   m_sin[494]  =  13'b1110011001001;     //494pi/512
   m_cos[494]  =  13'b1100010101101;     //494pi/512
   m_sin[495]  =  13'b1110011010011;     //495pi/512
   m_cos[495]  =  13'b1100010101000;     //495pi/512
   m_sin[496]  =  13'b1110011011110;     //496pi/512
   m_cos[496]  =  13'b1100010100100;     //496pi/512
   m_sin[497]  =  13'b1110011101000;     //497pi/512
   m_cos[497]  =  13'b1100010011111;     //497pi/512
   m_sin[498]  =  13'b1110011110011;     //498pi/512
   m_cos[498]  =  13'b1100010011011;     //498pi/512
   m_sin[499]  =  13'b1110011111101;     //499pi/512
   m_cos[499]  =  13'b1100010010111;     //499pi/512
   m_sin[500]  =  13'b1110100001000;     //500pi/512
   m_cos[500]  =  13'b1100010010010;     //500pi/512
   m_sin[501]  =  13'b1110100010010;     //501pi/512
   m_cos[501]  =  13'b1100010001110;     //501pi/512
   m_sin[502]  =  13'b1110100011101;     //502pi/512
   m_cos[502]  =  13'b1100010001010;     //502pi/512
   m_sin[503]  =  13'b1110100100111;     //503pi/512
   m_cos[503]  =  13'b1100010000110;     //503pi/512
   m_sin[504]  =  13'b1110100110010;     //504pi/512
   m_cos[504]  =  13'b1100010000010;     //504pi/512
   m_sin[505]  =  13'b1110100111100;     //505pi/512
   m_cos[505]  =  13'b1100001111110;     //505pi/512
   m_sin[506]  =  13'b1110101000111;     //506pi/512
   m_cos[506]  =  13'b1100001111010;     //506pi/512
   m_sin[507]  =  13'b1110101010010;     //507pi/512
   m_cos[507]  =  13'b1100001110110;     //507pi/512
   m_sin[508]  =  13'b1110101011100;     //508pi/512
   m_cos[508]  =  13'b1100001110011;     //508pi/512
   m_sin[509]  =  13'b1110101100111;     //509pi/512
   m_cos[509]  =  13'b1100001101111;     //509pi/512
   m_sin[510]  =  13'b1110101110010;     //510pi/512
   m_cos[510]  =  13'b1100001101011;     //510pi/512
   m_sin[511]  =  13'b1110101111100;     //511pi/512
   m_cos[511]  =  13'b1100001101000;     //511pi/512
end
endmodule
