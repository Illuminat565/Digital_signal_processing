module  M_TWIDLE_14_bit #(parameter SIZE =10) (
    input            en_modify, 
    input   [10:0]   rd_ptr_angle,

    output  signed [13:0]   cos_data,
    output  signed [13:0]   sin_data
 );


wire signed [13:0]  cos  [511:0];
wire signed [13:0]  sin  [511:0];

wire signed [13:0]  cos2  [511:0];
wire signed [13:0]  sin2  [511:0];

assign cos_data =   en_modify? cos2 [rd_ptr_angle] : cos [rd_ptr_angle];
assign sin_data =   en_modify? sin2 [rd_ptr_angle] : sin [rd_ptr_angle];

  assign sin[0]  =  14'b00000000000000;     //0pi/512
  assign cos[0]  =  14'b01000000000000;     //0pi/512
  assign sin[1]  =  14'b11111111100111;     //1pi/512
  assign cos[1]  =  14'b00111111111111;     //1pi/512
  assign sin[2]  =  14'b11111111001110;     //2pi/512
  assign cos[2]  =  14'b00111111111111;     //2pi/512
  assign sin[3]  =  14'b11111110110101;     //3pi/512
  assign cos[3]  =  14'b00111111111111;     //3pi/512
  assign sin[4]  =  14'b11111110011011;     //4pi/512
  assign cos[4]  =  14'b00111111111110;     //4pi/512
  assign sin[5]  =  14'b11111110000010;     //5pi/512
  assign cos[5]  =  14'b00111111111110;     //5pi/512
  assign sin[6]  =  14'b11111101101001;     //6pi/512
  assign cos[6]  =  14'b00111111111101;     //6pi/512
  assign sin[7]  =  14'b11111101010000;     //7pi/512
  assign cos[7]  =  14'b00111111111100;     //7pi/512
  assign sin[8]  =  14'b11111100110111;     //8pi/512
  assign cos[8]  =  14'b00111111111011;     //8pi/512
  assign sin[9]  =  14'b11111100011110;     //9pi/512
  assign cos[9]  =  14'b00111111111001;     //9pi/512
  assign sin[10]  =  14'b11111100000101;     //10pi/512
  assign cos[10]  =  14'b00111111111000;     //10pi/512
  assign sin[11]  =  14'b11111011101100;     //11pi/512
  assign cos[11]  =  14'b00111111110110;     //11pi/512
  assign sin[12]  =  14'b11111011010011;     //12pi/512
  assign cos[12]  =  14'b00111111110100;     //12pi/512
  assign sin[13]  =  14'b11111010111010;     //13pi/512
  assign cos[13]  =  14'b00111111110010;     //13pi/512
  assign sin[14]  =  14'b11111010100001;     //14pi/512
  assign cos[14]  =  14'b00111111110000;     //14pi/512
  assign sin[15]  =  14'b11111010001000;     //15pi/512
  assign cos[15]  =  14'b00111111101110;     //15pi/512
  assign sin[16]  =  14'b11111001101111;     //16pi/512
  assign cos[16]  =  14'b00111111101100;     //16pi/512
  assign sin[17]  =  14'b11111001010110;     //17pi/512
  assign cos[17]  =  14'b00111111101001;     //17pi/512
  assign sin[18]  =  14'b11111000111101;     //18pi/512
  assign cos[18]  =  14'b00111111100111;     //18pi/512
  assign sin[19]  =  14'b11111000100100;     //19pi/512
  assign cos[19]  =  14'b00111111100100;     //19pi/512
  assign sin[20]  =  14'b11111000001011;     //20pi/512
  assign cos[20]  =  14'b00111111100001;     //20pi/512
  assign sin[21]  =  14'b11110111110010;     //21pi/512
  assign cos[21]  =  14'b00111111011110;     //21pi/512
  assign sin[22]  =  14'b11110111011001;     //22pi/512
  assign cos[22]  =  14'b00111111011010;     //22pi/512
  assign sin[23]  =  14'b11110111000000;     //23pi/512
  assign cos[23]  =  14'b00111111010111;     //23pi/512
  assign sin[24]  =  14'b11110110100111;     //24pi/512
  assign cos[24]  =  14'b00111111010011;     //24pi/512
  assign sin[25]  =  14'b11110110001110;     //25pi/512
  assign cos[25]  =  14'b00111111001111;     //25pi/512
  assign sin[26]  =  14'b11110101110101;     //26pi/512
  assign cos[26]  =  14'b00111111001011;     //26pi/512
  assign sin[27]  =  14'b11110101011101;     //27pi/512
  assign cos[27]  =  14'b00111111000111;     //27pi/512
  assign sin[28]  =  14'b11110101000100;     //28pi/512
  assign cos[28]  =  14'b00111111000011;     //28pi/512
  assign sin[29]  =  14'b11110100101011;     //29pi/512
  assign cos[29]  =  14'b00111110111111;     //29pi/512
  assign sin[30]  =  14'b11110100010010;     //30pi/512
  assign cos[30]  =  14'b00111110111010;     //30pi/512
  assign sin[31]  =  14'b11110011111010;     //31pi/512
  assign cos[31]  =  14'b00111110110110;     //31pi/512
  assign sin[32]  =  14'b11110011100001;     //32pi/512
  assign cos[32]  =  14'b00111110110001;     //32pi/512
  assign sin[33]  =  14'b11110011001000;     //33pi/512
  assign cos[33]  =  14'b00111110101100;     //33pi/512
  assign sin[34]  =  14'b11110010110000;     //34pi/512
  assign cos[34]  =  14'b00111110100111;     //34pi/512
  assign sin[35]  =  14'b11110010010111;     //35pi/512
  assign cos[35]  =  14'b00111110100001;     //35pi/512
  assign sin[36]  =  14'b11110001111111;     //36pi/512
  assign cos[36]  =  14'b00111110011100;     //36pi/512
  assign sin[37]  =  14'b11110001100110;     //37pi/512
  assign cos[37]  =  14'b00111110010110;     //37pi/512
  assign sin[38]  =  14'b11110001001110;     //38pi/512
  assign cos[38]  =  14'b00111110010001;     //38pi/512
  assign sin[39]  =  14'b11110000110101;     //39pi/512
  assign cos[39]  =  14'b00111110001011;     //39pi/512
  assign sin[40]  =  14'b11110000011101;     //40pi/512
  assign cos[40]  =  14'b00111110000101;     //40pi/512
  assign sin[41]  =  14'b11110000000100;     //41pi/512
  assign cos[41]  =  14'b00111101111111;     //41pi/512
  assign sin[42]  =  14'b11101111101100;     //42pi/512
  assign cos[42]  =  14'b00111101111000;     //42pi/512
  assign sin[43]  =  14'b11101111010100;     //43pi/512
  assign cos[43]  =  14'b00111101110010;     //43pi/512
  assign sin[44]  =  14'b11101110111100;     //44pi/512
  assign cos[44]  =  14'b00111101101011;     //44pi/512
  assign sin[45]  =  14'b11101110100011;     //45pi/512
  assign cos[45]  =  14'b00111101100100;     //45pi/512
  assign sin[46]  =  14'b11101110001011;     //46pi/512
  assign cos[46]  =  14'b00111101011101;     //46pi/512
  assign sin[47]  =  14'b11101101110011;     //47pi/512
  assign cos[47]  =  14'b00111101010110;     //47pi/512
  assign sin[48]  =  14'b11101101011011;     //48pi/512
  assign cos[48]  =  14'b00111101001111;     //48pi/512
  assign sin[49]  =  14'b11101101000011;     //49pi/512
  assign cos[49]  =  14'b00111101001000;     //49pi/512
  assign sin[50]  =  14'b11101100101011;     //50pi/512
  assign cos[50]  =  14'b00111101000000;     //50pi/512
  assign sin[51]  =  14'b11101100010011;     //51pi/512
  assign cos[51]  =  14'b00111100111001;     //51pi/512
  assign sin[52]  =  14'b11101011111011;     //52pi/512
  assign cos[52]  =  14'b00111100110001;     //52pi/512
  assign sin[53]  =  14'b11101011100011;     //53pi/512
  assign cos[53]  =  14'b00111100101001;     //53pi/512
  assign sin[54]  =  14'b11101011001100;     //54pi/512
  assign cos[54]  =  14'b00111100100001;     //54pi/512
  assign sin[55]  =  14'b11101010110100;     //55pi/512
  assign cos[55]  =  14'b00111100011000;     //55pi/512
  assign sin[56]  =  14'b11101010011100;     //56pi/512
  assign cos[56]  =  14'b00111100010000;     //56pi/512
  assign sin[57]  =  14'b11101010000100;     //57pi/512
  assign cos[57]  =  14'b00111100001000;     //57pi/512
  assign sin[58]  =  14'b11101001101101;     //58pi/512
  assign cos[58]  =  14'b00111011111111;     //58pi/512
  assign sin[59]  =  14'b11101001010101;     //59pi/512
  assign cos[59]  =  14'b00111011110110;     //59pi/512
  assign sin[60]  =  14'b11101000111110;     //60pi/512
  assign cos[60]  =  14'b00111011101101;     //60pi/512
  assign sin[61]  =  14'b11101000100110;     //61pi/512
  assign cos[61]  =  14'b00111011100100;     //61pi/512
  assign sin[62]  =  14'b11101000001111;     //62pi/512
  assign cos[62]  =  14'b00111011011011;     //62pi/512
  assign sin[63]  =  14'b11100111111000;     //63pi/512
  assign cos[63]  =  14'b00111011010001;     //63pi/512
  assign sin[64]  =  14'b11100111100001;     //64pi/512
  assign cos[64]  =  14'b00111011001000;     //64pi/512
  assign sin[65]  =  14'b11100111001001;     //65pi/512
  assign cos[65]  =  14'b00111010111110;     //65pi/512
  assign sin[66]  =  14'b11100110110010;     //66pi/512
  assign cos[66]  =  14'b00111010110100;     //66pi/512
  assign sin[67]  =  14'b11100110011011;     //67pi/512
  assign cos[67]  =  14'b00111010101010;     //67pi/512
  assign sin[68]  =  14'b11100110000100;     //68pi/512
  assign cos[68]  =  14'b00111010100000;     //68pi/512
  assign sin[69]  =  14'b11100101101101;     //69pi/512
  assign cos[69]  =  14'b00111010010110;     //69pi/512
  assign sin[70]  =  14'b11100101010110;     //70pi/512
  assign cos[70]  =  14'b00111010001011;     //70pi/512
  assign sin[71]  =  14'b11100100111111;     //71pi/512
  assign cos[71]  =  14'b00111010000001;     //71pi/512
  assign sin[72]  =  14'b11100100101001;     //72pi/512
  assign cos[72]  =  14'b00111001110110;     //72pi/512
  assign sin[73]  =  14'b11100100010010;     //73pi/512
  assign cos[73]  =  14'b00111001101011;     //73pi/512
  assign sin[74]  =  14'b11100011111011;     //74pi/512
  assign cos[74]  =  14'b00111001100000;     //74pi/512
  assign sin[75]  =  14'b11100011100101;     //75pi/512
  assign cos[75]  =  14'b00111001010101;     //75pi/512
  assign sin[76]  =  14'b11100011001110;     //76pi/512
  assign cos[76]  =  14'b00111001001010;     //76pi/512
  assign sin[77]  =  14'b11100010111000;     //77pi/512
  assign cos[77]  =  14'b00111000111111;     //77pi/512
  assign sin[78]  =  14'b11100010100010;     //78pi/512
  assign cos[78]  =  14'b00111000110011;     //78pi/512
  assign sin[79]  =  14'b11100010001011;     //79pi/512
  assign cos[79]  =  14'b00111000101000;     //79pi/512
  assign sin[80]  =  14'b11100001110101;     //80pi/512
  assign cos[80]  =  14'b00111000011100;     //80pi/512
  assign sin[81]  =  14'b11100001011111;     //81pi/512
  assign cos[81]  =  14'b00111000010000;     //81pi/512
  assign sin[82]  =  14'b11100001001001;     //82pi/512
  assign cos[82]  =  14'b00111000000100;     //82pi/512
  assign sin[83]  =  14'b11100000110011;     //83pi/512
  assign cos[83]  =  14'b00110111111000;     //83pi/512
  assign sin[84]  =  14'b11100000011101;     //84pi/512
  assign cos[84]  =  14'b00110111101011;     //84pi/512
  assign sin[85]  =  14'b11100000000111;     //85pi/512
  assign cos[85]  =  14'b00110111011111;     //85pi/512
  assign sin[86]  =  14'b11011111110010;     //86pi/512
  assign cos[86]  =  14'b00110111010010;     //86pi/512
  assign sin[87]  =  14'b11011111011100;     //87pi/512
  assign cos[87]  =  14'b00110111000110;     //87pi/512
  assign sin[88]  =  14'b11011111000110;     //88pi/512
  assign cos[88]  =  14'b00110110111001;     //88pi/512
  assign sin[89]  =  14'b11011110110001;     //89pi/512
  assign cos[89]  =  14'b00110110101100;     //89pi/512
  assign sin[90]  =  14'b11011110011011;     //90pi/512
  assign cos[90]  =  14'b00110110011111;     //90pi/512
  assign sin[91]  =  14'b11011110000110;     //91pi/512
  assign cos[91]  =  14'b00110110010001;     //91pi/512
  assign sin[92]  =  14'b11011101110001;     //92pi/512
  assign cos[92]  =  14'b00110110000100;     //92pi/512
  assign sin[93]  =  14'b11011101011011;     //93pi/512
  assign cos[93]  =  14'b00110101110111;     //93pi/512
  assign sin[94]  =  14'b11011101000110;     //94pi/512
  assign cos[94]  =  14'b00110101101001;     //94pi/512
  assign sin[95]  =  14'b11011100110001;     //95pi/512
  assign cos[95]  =  14'b00110101011011;     //95pi/512
  assign sin[96]  =  14'b11011100011100;     //96pi/512
  assign cos[96]  =  14'b00110101001101;     //96pi/512
  assign sin[97]  =  14'b11011100001000;     //97pi/512
  assign cos[97]  =  14'b00110100111111;     //97pi/512
  assign sin[98]  =  14'b11011011110011;     //98pi/512
  assign cos[98]  =  14'b00110100110001;     //98pi/512
  assign sin[99]  =  14'b11011011011110;     //99pi/512
  assign cos[99]  =  14'b00110100100011;     //99pi/512
  assign sin[100]  =  14'b11011011001001;     //100pi/512
  assign cos[100]  =  14'b00110100010100;     //100pi/512
  assign sin[101]  =  14'b11011010110101;     //101pi/512
  assign cos[101]  =  14'b00110100000110;     //101pi/512
  assign sin[102]  =  14'b11011010100001;     //102pi/512
  assign cos[102]  =  14'b00110011110111;     //102pi/512
  assign sin[103]  =  14'b11011010001100;     //103pi/512
  assign cos[103]  =  14'b00110011101000;     //103pi/512
  assign sin[104]  =  14'b11011001111000;     //104pi/512
  assign cos[104]  =  14'b00110011011001;     //104pi/512
  assign sin[105]  =  14'b11011001100100;     //105pi/512
  assign cos[105]  =  14'b00110011001010;     //105pi/512
  assign sin[106]  =  14'b11011001010000;     //106pi/512
  assign cos[106]  =  14'b00110010111011;     //106pi/512
  assign sin[107]  =  14'b11011000111100;     //107pi/512
  assign cos[107]  =  14'b00110010101100;     //107pi/512
  assign sin[108]  =  14'b11011000101000;     //108pi/512
  assign cos[108]  =  14'b00110010011101;     //108pi/512
  assign sin[109]  =  14'b11011000010100;     //109pi/512
  assign cos[109]  =  14'b00110010001101;     //109pi/512
  assign sin[110]  =  14'b11011000000001;     //110pi/512
  assign cos[110]  =  14'b00110001111101;     //110pi/512
  assign sin[111]  =  14'b11010111101101;     //111pi/512
  assign cos[111]  =  14'b00110001101110;     //111pi/512
  assign sin[112]  =  14'b11010111011010;     //112pi/512
  assign cos[112]  =  14'b00110001011110;     //112pi/512
  assign sin[113]  =  14'b11010111000110;     //113pi/512
  assign cos[113]  =  14'b00110001001110;     //113pi/512
  assign sin[114]  =  14'b11010110110011;     //114pi/512
  assign cos[114]  =  14'b00110000111110;     //114pi/512
  assign sin[115]  =  14'b11010110100000;     //115pi/512
  assign cos[115]  =  14'b00110000101101;     //115pi/512
  assign sin[116]  =  14'b11010110001101;     //116pi/512
  assign cos[116]  =  14'b00110000011101;     //116pi/512
  assign sin[117]  =  14'b11010101111010;     //117pi/512
  assign cos[117]  =  14'b00110000001101;     //117pi/512
  assign sin[118]  =  14'b11010101100111;     //118pi/512
  assign cos[118]  =  14'b00101111111100;     //118pi/512
  assign sin[119]  =  14'b11010101010100;     //119pi/512
  assign cos[119]  =  14'b00101111101011;     //119pi/512
  assign sin[120]  =  14'b11010101000001;     //120pi/512
  assign cos[120]  =  14'b00101111011010;     //120pi/512
  assign sin[121]  =  14'b11010100101111;     //121pi/512
  assign cos[121]  =  14'b00101111001010;     //121pi/512
  assign sin[122]  =  14'b11010100011100;     //122pi/512
  assign cos[122]  =  14'b00101110111000;     //122pi/512
  assign sin[123]  =  14'b11010100001010;     //123pi/512
  assign cos[123]  =  14'b00101110100111;     //123pi/512
  assign sin[124]  =  14'b11010011111000;     //124pi/512
  assign cos[124]  =  14'b00101110010110;     //124pi/512
  assign sin[125]  =  14'b11010011100101;     //125pi/512
  assign cos[125]  =  14'b00101110000101;     //125pi/512
  assign sin[126]  =  14'b11010011010011;     //126pi/512
  assign cos[126]  =  14'b00101101110011;     //126pi/512
  assign sin[127]  =  14'b11010011000010;     //127pi/512
  assign cos[127]  =  14'b00101101100010;     //127pi/512
  assign sin[128]  =  14'b11010010110000;     //128pi/512
  assign cos[128]  =  14'b00101101010000;     //128pi/512
  assign sin[129]  =  14'b11010010011110;     //129pi/512
  assign cos[129]  =  14'b00101100111110;     //129pi/512
  assign sin[130]  =  14'b11010010001100;     //130pi/512
  assign cos[130]  =  14'b00101100101100;     //130pi/512
  assign sin[131]  =  14'b11010001111011;     //131pi/512
  assign cos[131]  =  14'b00101100011010;     //131pi/512
  assign sin[132]  =  14'b11010001101001;     //132pi/512
  assign cos[132]  =  14'b00101100001000;     //132pi/512
  assign sin[133]  =  14'b11010001011000;     //133pi/512
  assign cos[133]  =  14'b00101011110110;     //133pi/512
  assign sin[134]  =  14'b11010001000111;     //134pi/512
  assign cos[134]  =  14'b00101011100011;     //134pi/512
  assign sin[135]  =  14'b11010000110110;     //135pi/512
  assign cos[135]  =  14'b00101011010001;     //135pi/512
  assign sin[136]  =  14'b11010000100101;     //136pi/512
  assign cos[136]  =  14'b00101010111110;     //136pi/512
  assign sin[137]  =  14'b11010000010100;     //137pi/512
  assign cos[137]  =  14'b00101010101100;     //137pi/512
  assign sin[138]  =  14'b11010000000100;     //138pi/512
  assign cos[138]  =  14'b00101010011001;     //138pi/512
  assign sin[139]  =  14'b11001111110011;     //139pi/512
  assign cos[139]  =  14'b00101010000110;     //139pi/512
  assign sin[140]  =  14'b11001111100010;     //140pi/512
  assign cos[140]  =  14'b00101001110011;     //140pi/512
  assign sin[141]  =  14'b11001111010010;     //141pi/512
  assign cos[141]  =  14'b00101001100000;     //141pi/512
  assign sin[142]  =  14'b11001111000010;     //142pi/512
  assign cos[142]  =  14'b00101001001101;     //142pi/512
  assign sin[143]  =  14'b11001110110010;     //143pi/512
  assign cos[143]  =  14'b00101000111001;     //143pi/512
  assign sin[144]  =  14'b11001110100010;     //144pi/512
  assign cos[144]  =  14'b00101000100110;     //144pi/512
  assign sin[145]  =  14'b11001110010010;     //145pi/512
  assign cos[145]  =  14'b00101000010010;     //145pi/512
  assign sin[146]  =  14'b11001110000010;     //146pi/512
  assign cos[146]  =  14'b00100111111111;     //146pi/512
  assign sin[147]  =  14'b11001101110010;     //147pi/512
  assign cos[147]  =  14'b00100111101011;     //147pi/512
  assign sin[148]  =  14'b11001101100011;     //148pi/512
  assign cos[148]  =  14'b00100111010111;     //148pi/512
  assign sin[149]  =  14'b11001101010100;     //149pi/512
  assign cos[149]  =  14'b00100111000100;     //149pi/512
  assign sin[150]  =  14'b11001101000100;     //150pi/512
  assign cos[150]  =  14'b00100110110000;     //150pi/512
  assign sin[151]  =  14'b11001100110101;     //151pi/512
  assign cos[151]  =  14'b00100110011100;     //151pi/512
  assign sin[152]  =  14'b11001100100110;     //152pi/512
  assign cos[152]  =  14'b00100110000111;     //152pi/512
  assign sin[153]  =  14'b11001100010111;     //153pi/512
  assign cos[153]  =  14'b00100101110011;     //153pi/512
  assign sin[154]  =  14'b11001100001000;     //154pi/512
  assign cos[154]  =  14'b00100101011111;     //154pi/512
  assign sin[155]  =  14'b11001011111010;     //155pi/512
  assign cos[155]  =  14'b00100101001011;     //155pi/512
  assign sin[156]  =  14'b11001011101011;     //156pi/512
  assign cos[156]  =  14'b00100100110110;     //156pi/512
  assign sin[157]  =  14'b11001011011101;     //157pi/512
  assign cos[157]  =  14'b00100100100001;     //157pi/512
  assign sin[158]  =  14'b11001011001110;     //158pi/512
  assign cos[158]  =  14'b00100100001101;     //158pi/512
  assign sin[159]  =  14'b11001011000000;     //159pi/512
  assign cos[159]  =  14'b00100011111000;     //159pi/512
  assign sin[160]  =  14'b11001010110010;     //160pi/512
  assign cos[160]  =  14'b00100011100011;     //160pi/512
  assign sin[161]  =  14'b11001010100100;     //161pi/512
  assign cos[161]  =  14'b00100011001110;     //161pi/512
  assign sin[162]  =  14'b11001010010111;     //162pi/512
  assign cos[162]  =  14'b00100010111001;     //162pi/512
  assign sin[163]  =  14'b11001010001001;     //163pi/512
  assign cos[163]  =  14'b00100010100100;     //163pi/512
  assign sin[164]  =  14'b11001001111011;     //164pi/512
  assign cos[164]  =  14'b00100010001111;     //164pi/512
  assign sin[165]  =  14'b11001001101110;     //165pi/512
  assign cos[165]  =  14'b00100001111010;     //165pi/512
  assign sin[166]  =  14'b11001001100001;     //166pi/512
  assign cos[166]  =  14'b00100001100100;     //166pi/512
  assign sin[167]  =  14'b11001001010100;     //167pi/512
  assign cos[167]  =  14'b00100001001111;     //167pi/512
  assign sin[168]  =  14'b11001001000111;     //168pi/512
  assign cos[168]  =  14'b00100000111001;     //168pi/512
  assign sin[169]  =  14'b11001000111010;     //169pi/512
  assign cos[169]  =  14'b00100000100100;     //169pi/512
  assign sin[170]  =  14'b11001000101101;     //170pi/512
  assign cos[170]  =  14'b00100000001110;     //170pi/512
  assign sin[171]  =  14'b11001000100001;     //171pi/512
  assign cos[171]  =  14'b00011111111000;     //171pi/512
  assign sin[172]  =  14'b11001000010100;     //172pi/512
  assign cos[172]  =  14'b00011111100010;     //172pi/512
  assign sin[173]  =  14'b11001000001000;     //173pi/512
  assign cos[173]  =  14'b00011111001101;     //173pi/512
  assign sin[174]  =  14'b11000111111100;     //174pi/512
  assign cos[174]  =  14'b00011110110111;     //174pi/512
  assign sin[175]  =  14'b11000111110000;     //175pi/512
  assign cos[175]  =  14'b00011110100000;     //175pi/512
  assign sin[176]  =  14'b11000111100100;     //176pi/512
  assign cos[176]  =  14'b00011110001010;     //176pi/512
  assign sin[177]  =  14'b11000111011000;     //177pi/512
  assign cos[177]  =  14'b00011101110100;     //177pi/512
  assign sin[178]  =  14'b11000111001100;     //178pi/512
  assign cos[178]  =  14'b00011101011110;     //178pi/512
  assign sin[179]  =  14'b11000111000001;     //179pi/512
  assign cos[179]  =  14'b00011101001000;     //179pi/512
  assign sin[180]  =  14'b11000110110101;     //180pi/512
  assign cos[180]  =  14'b00011100110001;     //180pi/512
  assign sin[181]  =  14'b11000110101010;     //181pi/512
  assign cos[181]  =  14'b00011100011011;     //181pi/512
  assign sin[182]  =  14'b11000110011111;     //182pi/512
  assign cos[182]  =  14'b00011100000100;     //182pi/512
  assign sin[183]  =  14'b11000110010100;     //183pi/512
  assign cos[183]  =  14'b00011011101101;     //183pi/512
  assign sin[184]  =  14'b11000110001001;     //184pi/512
  assign cos[184]  =  14'b00011011010111;     //184pi/512
  assign sin[185]  =  14'b11000101111111;     //185pi/512
  assign cos[185]  =  14'b00011011000000;     //185pi/512
  assign sin[186]  =  14'b11000101110100;     //186pi/512
  assign cos[186]  =  14'b00011010101001;     //186pi/512
  assign sin[187]  =  14'b11000101101010;     //187pi/512
  assign cos[187]  =  14'b00011010010010;     //187pi/512
  assign sin[188]  =  14'b11000101011111;     //188pi/512
  assign cos[188]  =  14'b00011001111011;     //188pi/512
  assign sin[189]  =  14'b11000101010101;     //189pi/512
  assign cos[189]  =  14'b00011001100100;     //189pi/512
  assign sin[190]  =  14'b11000101001011;     //190pi/512
  assign cos[190]  =  14'b00011001001101;     //190pi/512
  assign sin[191]  =  14'b11000101000001;     //191pi/512
  assign cos[191]  =  14'b00011000110110;     //191pi/512
  assign sin[192]  =  14'b11000100111000;     //192pi/512
  assign cos[192]  =  14'b00011000011111;     //192pi/512
  assign sin[193]  =  14'b11000100101110;     //193pi/512
  assign cos[193]  =  14'b00011000001000;     //193pi/512
  assign sin[194]  =  14'b11000100100101;     //194pi/512
  assign cos[194]  =  14'b00010111110000;     //194pi/512
  assign sin[195]  =  14'b11000100011100;     //195pi/512
  assign cos[195]  =  14'b00010111011001;     //195pi/512
  assign sin[196]  =  14'b11000100010010;     //196pi/512
  assign cos[196]  =  14'b00010111000010;     //196pi/512
  assign sin[197]  =  14'b11000100001001;     //197pi/512
  assign cos[197]  =  14'b00010110101010;     //197pi/512
  assign sin[198]  =  14'b11000100000001;     //198pi/512
  assign cos[198]  =  14'b00010110010011;     //198pi/512
  assign sin[199]  =  14'b11000011111000;     //199pi/512
  assign cos[199]  =  14'b00010101111011;     //199pi/512
  assign sin[200]  =  14'b11000011101111;     //200pi/512
  assign cos[200]  =  14'b00010101100011;     //200pi/512
  assign sin[201]  =  14'b11000011100111;     //201pi/512
  assign cos[201]  =  14'b00010101001100;     //201pi/512
  assign sin[202]  =  14'b11000011011111;     //202pi/512
  assign cos[202]  =  14'b00010100110100;     //202pi/512
  assign sin[203]  =  14'b11000011010111;     //203pi/512
  assign cos[203]  =  14'b00010100011100;     //203pi/512
  assign sin[204]  =  14'b11000011001111;     //204pi/512
  assign cos[204]  =  14'b00010100000100;     //204pi/512
  assign sin[205]  =  14'b11000011000111;     //205pi/512
  assign cos[205]  =  14'b00010011101100;     //205pi/512
  assign sin[206]  =  14'b11000010111111;     //206pi/512
  assign cos[206]  =  14'b00010011010101;     //206pi/512
  assign sin[207]  =  14'b11000010111000;     //207pi/512
  assign cos[207]  =  14'b00010010111101;     //207pi/512
  assign sin[208]  =  14'b11000010110000;     //208pi/512
  assign cos[208]  =  14'b00010010100101;     //208pi/512
  assign sin[209]  =  14'b11000010101001;     //209pi/512
  assign cos[209]  =  14'b00010010001100;     //209pi/512
  assign sin[210]  =  14'b11000010100010;     //210pi/512
  assign cos[210]  =  14'b00010001110100;     //210pi/512
  assign sin[211]  =  14'b11000010011011;     //211pi/512
  assign cos[211]  =  14'b00010001011100;     //211pi/512
  assign sin[212]  =  14'b11000010010100;     //212pi/512
  assign cos[212]  =  14'b00010001000100;     //212pi/512
  assign sin[213]  =  14'b11000010001110;     //213pi/512
  assign cos[213]  =  14'b00010000101100;     //213pi/512
  assign sin[214]  =  14'b11000010000111;     //214pi/512
  assign cos[214]  =  14'b00010000010011;     //214pi/512
  assign sin[215]  =  14'b11000010000001;     //215pi/512
  assign cos[215]  =  14'b00001111111011;     //215pi/512
  assign sin[216]  =  14'b11000001111011;     //216pi/512
  assign cos[216]  =  14'b00001111100011;     //216pi/512
  assign sin[217]  =  14'b11000001110101;     //217pi/512
  assign cos[217]  =  14'b00001111001010;     //217pi/512
  assign sin[218]  =  14'b11000001101111;     //218pi/512
  assign cos[218]  =  14'b00001110110010;     //218pi/512
  assign sin[219]  =  14'b11000001101001;     //219pi/512
  assign cos[219]  =  14'b00001110011001;     //219pi/512
  assign sin[220]  =  14'b11000001100100;     //220pi/512
  assign cos[220]  =  14'b00001110000001;     //220pi/512
  assign sin[221]  =  14'b11000001011110;     //221pi/512
  assign cos[221]  =  14'b00001101101000;     //221pi/512
  assign sin[222]  =  14'b11000001011001;     //222pi/512
  assign cos[222]  =  14'b00001101010000;     //222pi/512
  assign sin[223]  =  14'b11000001010100;     //223pi/512
  assign cos[223]  =  14'b00001100110111;     //223pi/512
  assign sin[224]  =  14'b11000001001111;     //224pi/512
  assign cos[224]  =  14'b00001100011111;     //224pi/512
  assign sin[225]  =  14'b11000001001010;     //225pi/512
  assign cos[225]  =  14'b00001100000110;     //225pi/512
  assign sin[226]  =  14'b11000001000101;     //226pi/512
  assign cos[226]  =  14'b00001011101101;     //226pi/512
  assign sin[227]  =  14'b11000001000001;     //227pi/512
  assign cos[227]  =  14'b00001011010101;     //227pi/512
  assign sin[228]  =  14'b11000000111100;     //228pi/512
  assign cos[228]  =  14'b00001010111100;     //228pi/512
  assign sin[229]  =  14'b11000000111000;     //229pi/512
  assign cos[229]  =  14'b00001010100011;     //229pi/512
  assign sin[230]  =  14'b11000000110100;     //230pi/512
  assign cos[230]  =  14'b00001010001010;     //230pi/512
  assign sin[231]  =  14'b11000000110000;     //231pi/512
  assign cos[231]  =  14'b00001001110001;     //231pi/512
  assign sin[232]  =  14'b11000000101100;     //232pi/512
  assign cos[232]  =  14'b00001001011001;     //232pi/512
  assign sin[233]  =  14'b11000000101001;     //233pi/512
  assign cos[233]  =  14'b00001001000000;     //233pi/512
  assign sin[234]  =  14'b11000000100101;     //234pi/512
  assign cos[234]  =  14'b00001000100111;     //234pi/512
  assign sin[235]  =  14'b11000000100010;     //235pi/512
  assign cos[235]  =  14'b00001000001110;     //235pi/512
  assign sin[236]  =  14'b11000000011111;     //236pi/512
  assign cos[236]  =  14'b00000111110101;     //236pi/512
  assign sin[237]  =  14'b11000000011100;     //237pi/512
  assign cos[237]  =  14'b00000111011100;     //237pi/512
  assign sin[238]  =  14'b11000000011001;     //238pi/512
  assign cos[238]  =  14'b00000111000011;     //238pi/512
  assign sin[239]  =  14'b11000000010110;     //239pi/512
  assign cos[239]  =  14'b00000110101010;     //239pi/512
  assign sin[240]  =  14'b11000000010100;     //240pi/512
  assign cos[240]  =  14'b00000110010001;     //240pi/512
  assign sin[241]  =  14'b11000000010001;     //241pi/512
  assign cos[241]  =  14'b00000101111000;     //241pi/512
  assign sin[242]  =  14'b11000000001111;     //242pi/512
  assign cos[242]  =  14'b00000101011111;     //242pi/512
  assign sin[243]  =  14'b11000000001101;     //243pi/512
  assign cos[243]  =  14'b00000101000110;     //243pi/512
  assign sin[244]  =  14'b11000000001011;     //244pi/512
  assign cos[244]  =  14'b00000100101101;     //244pi/512
  assign sin[245]  =  14'b11000000001001;     //245pi/512
  assign cos[245]  =  14'b00000100010100;     //245pi/512
  assign sin[246]  =  14'b11000000001000;     //246pi/512
  assign cos[246]  =  14'b00000011111011;     //246pi/512
  assign sin[247]  =  14'b11000000000110;     //247pi/512
  assign cos[247]  =  14'b00000011100010;     //247pi/512
  assign sin[248]  =  14'b11000000000101;     //248pi/512
  assign cos[248]  =  14'b00000011001000;     //248pi/512
  assign sin[249]  =  14'b11000000000100;     //249pi/512
  assign cos[249]  =  14'b00000010101111;     //249pi/512
  assign sin[250]  =  14'b11000000000011;     //250pi/512
  assign cos[250]  =  14'b00000010010110;     //250pi/512
  assign sin[251]  =  14'b11000000000010;     //251pi/512
  assign cos[251]  =  14'b00000001111101;     //251pi/512
  assign sin[252]  =  14'b11000000000001;     //252pi/512
  assign cos[252]  =  14'b00000001100100;     //252pi/512
  assign sin[253]  =  14'b11000000000001;     //253pi/512
  assign cos[253]  =  14'b00000001001011;     //253pi/512
  assign sin[254]  =  14'b11000000000000;     //254pi/512
  assign cos[254]  =  14'b00000000110010;     //254pi/512
  assign sin[255]  =  14'b11000000000000;     //255pi/512
  assign cos[255]  =  14'b00000000011001;     //255pi/512
  assign sin[256]  =  14'b11000000000000;     //256pi/512
  assign cos[256]  =  14'b00000000000000;     //256pi/512
  assign sin[257]  =  14'b11000000000000;     //257pi/512
  assign cos[257]  =  14'b11111111100111;     //257pi/512
  assign sin[258]  =  14'b11000000000000;     //258pi/512
  assign cos[258]  =  14'b11111111001110;     //258pi/512
  assign sin[259]  =  14'b11000000000001;     //259pi/512
  assign cos[259]  =  14'b11111110110101;     //259pi/512
  assign sin[260]  =  14'b11000000000001;     //260pi/512
  assign cos[260]  =  14'b11111110011011;     //260pi/512
  assign sin[261]  =  14'b11000000000010;     //261pi/512
  assign cos[261]  =  14'b11111110000010;     //261pi/512
  assign sin[262]  =  14'b11000000000011;     //262pi/512
  assign cos[262]  =  14'b11111101101001;     //262pi/512
  assign sin[263]  =  14'b11000000000100;     //263pi/512
  assign cos[263]  =  14'b11111101010000;     //263pi/512
  assign sin[264]  =  14'b11000000000101;     //264pi/512
  assign cos[264]  =  14'b11111100110111;     //264pi/512
  assign sin[265]  =  14'b11000000000110;     //265pi/512
  assign cos[265]  =  14'b11111100011110;     //265pi/512
  assign sin[266]  =  14'b11000000001000;     //266pi/512
  assign cos[266]  =  14'b11111100000101;     //266pi/512
  assign sin[267]  =  14'b11000000001001;     //267pi/512
  assign cos[267]  =  14'b11111011101100;     //267pi/512
  assign sin[268]  =  14'b11000000001011;     //268pi/512
  assign cos[268]  =  14'b11111011010011;     //268pi/512
  assign sin[269]  =  14'b11000000001101;     //269pi/512
  assign cos[269]  =  14'b11111010111010;     //269pi/512
  assign sin[270]  =  14'b11000000001111;     //270pi/512
  assign cos[270]  =  14'b11111010100001;     //270pi/512
  assign sin[271]  =  14'b11000000010001;     //271pi/512
  assign cos[271]  =  14'b11111010001000;     //271pi/512
  assign sin[272]  =  14'b11000000010100;     //272pi/512
  assign cos[272]  =  14'b11111001101111;     //272pi/512
  assign sin[273]  =  14'b11000000010110;     //273pi/512
  assign cos[273]  =  14'b11111001010110;     //273pi/512
  assign sin[274]  =  14'b11000000011001;     //274pi/512
  assign cos[274]  =  14'b11111000111101;     //274pi/512
  assign sin[275]  =  14'b11000000011100;     //275pi/512
  assign cos[275]  =  14'b11111000100100;     //275pi/512
  assign sin[276]  =  14'b11000000011111;     //276pi/512
  assign cos[276]  =  14'b11111000001011;     //276pi/512
  assign sin[277]  =  14'b11000000100010;     //277pi/512
  assign cos[277]  =  14'b11110111110010;     //277pi/512
  assign sin[278]  =  14'b11000000100101;     //278pi/512
  assign cos[278]  =  14'b11110111011001;     //278pi/512
  assign sin[279]  =  14'b11000000101001;     //279pi/512
  assign cos[279]  =  14'b11110111000000;     //279pi/512
  assign sin[280]  =  14'b11000000101100;     //280pi/512
  assign cos[280]  =  14'b11110110100111;     //280pi/512
  assign sin[281]  =  14'b11000000110000;     //281pi/512
  assign cos[281]  =  14'b11110110001110;     //281pi/512
  assign sin[282]  =  14'b11000000110100;     //282pi/512
  assign cos[282]  =  14'b11110101110101;     //282pi/512
  assign sin[283]  =  14'b11000000111000;     //283pi/512
  assign cos[283]  =  14'b11110101011101;     //283pi/512
  assign sin[284]  =  14'b11000000111100;     //284pi/512
  assign cos[284]  =  14'b11110101000100;     //284pi/512
  assign sin[285]  =  14'b11000001000001;     //285pi/512
  assign cos[285]  =  14'b11110100101011;     //285pi/512
  assign sin[286]  =  14'b11000001000101;     //286pi/512
  assign cos[286]  =  14'b11110100010010;     //286pi/512
  assign sin[287]  =  14'b11000001001010;     //287pi/512
  assign cos[287]  =  14'b11110011111010;     //287pi/512
  assign sin[288]  =  14'b11000001001111;     //288pi/512
  assign cos[288]  =  14'b11110011100001;     //288pi/512
  assign sin[289]  =  14'b11000001010100;     //289pi/512
  assign cos[289]  =  14'b11110011001000;     //289pi/512
  assign sin[290]  =  14'b11000001011001;     //290pi/512
  assign cos[290]  =  14'b11110010110000;     //290pi/512
  assign sin[291]  =  14'b11000001011110;     //291pi/512
  assign cos[291]  =  14'b11110010010111;     //291pi/512
  assign sin[292]  =  14'b11000001100100;     //292pi/512
  assign cos[292]  =  14'b11110001111111;     //292pi/512
  assign sin[293]  =  14'b11000001101001;     //293pi/512
  assign cos[293]  =  14'b11110001100110;     //293pi/512
  assign sin[294]  =  14'b11000001101111;     //294pi/512
  assign cos[294]  =  14'b11110001001110;     //294pi/512
  assign sin[295]  =  14'b11000001110101;     //295pi/512
  assign cos[295]  =  14'b11110000110101;     //295pi/512
  assign sin[296]  =  14'b11000001111011;     //296pi/512
  assign cos[296]  =  14'b11110000011101;     //296pi/512
  assign sin[297]  =  14'b11000010000001;     //297pi/512
  assign cos[297]  =  14'b11110000000100;     //297pi/512
  assign sin[298]  =  14'b11000010000111;     //298pi/512
  assign cos[298]  =  14'b11101111101100;     //298pi/512
  assign sin[299]  =  14'b11000010001110;     //299pi/512
  assign cos[299]  =  14'b11101111010100;     //299pi/512
  assign sin[300]  =  14'b11000010010100;     //300pi/512
  assign cos[300]  =  14'b11101110111100;     //300pi/512
  assign sin[301]  =  14'b11000010011011;     //301pi/512
  assign cos[301]  =  14'b11101110100011;     //301pi/512
  assign sin[302]  =  14'b11000010100010;     //302pi/512
  assign cos[302]  =  14'b11101110001011;     //302pi/512
  assign sin[303]  =  14'b11000010101001;     //303pi/512
  assign cos[303]  =  14'b11101101110011;     //303pi/512
  assign sin[304]  =  14'b11000010110000;     //304pi/512
  assign cos[304]  =  14'b11101101011011;     //304pi/512
  assign sin[305]  =  14'b11000010111000;     //305pi/512
  assign cos[305]  =  14'b11101101000011;     //305pi/512
  assign sin[306]  =  14'b11000010111111;     //306pi/512
  assign cos[306]  =  14'b11101100101011;     //306pi/512
  assign sin[307]  =  14'b11000011000111;     //307pi/512
  assign cos[307]  =  14'b11101100010011;     //307pi/512
  assign sin[308]  =  14'b11000011001111;     //308pi/512
  assign cos[308]  =  14'b11101011111011;     //308pi/512
  assign sin[309]  =  14'b11000011010111;     //309pi/512
  assign cos[309]  =  14'b11101011100011;     //309pi/512
  assign sin[310]  =  14'b11000011011111;     //310pi/512
  assign cos[310]  =  14'b11101011001100;     //310pi/512
  assign sin[311]  =  14'b11000011100111;     //311pi/512
  assign cos[311]  =  14'b11101010110100;     //311pi/512
  assign sin[312]  =  14'b11000011101111;     //312pi/512
  assign cos[312]  =  14'b11101010011100;     //312pi/512
  assign sin[313]  =  14'b11000011111000;     //313pi/512
  assign cos[313]  =  14'b11101010000100;     //313pi/512
  assign sin[314]  =  14'b11000100000001;     //314pi/512
  assign cos[314]  =  14'b11101001101101;     //314pi/512
  assign sin[315]  =  14'b11000100001001;     //315pi/512
  assign cos[315]  =  14'b11101001010101;     //315pi/512
  assign sin[316]  =  14'b11000100010010;     //316pi/512
  assign cos[316]  =  14'b11101000111110;     //316pi/512
  assign sin[317]  =  14'b11000100011100;     //317pi/512
  assign cos[317]  =  14'b11101000100110;     //317pi/512
  assign sin[318]  =  14'b11000100100101;     //318pi/512
  assign cos[318]  =  14'b11101000001111;     //318pi/512
  assign sin[319]  =  14'b11000100101110;     //319pi/512
  assign cos[319]  =  14'b11100111111000;     //319pi/512
  assign sin[320]  =  14'b11000100111000;     //320pi/512
  assign cos[320]  =  14'b11100111100001;     //320pi/512
  assign sin[321]  =  14'b11000101000001;     //321pi/512
  assign cos[321]  =  14'b11100111001001;     //321pi/512
  assign sin[322]  =  14'b11000101001011;     //322pi/512
  assign cos[322]  =  14'b11100110110010;     //322pi/512
  assign sin[323]  =  14'b11000101010101;     //323pi/512
  assign cos[323]  =  14'b11100110011011;     //323pi/512
  assign sin[324]  =  14'b11000101011111;     //324pi/512
  assign cos[324]  =  14'b11100110000100;     //324pi/512
  assign sin[325]  =  14'b11000101101010;     //325pi/512
  assign cos[325]  =  14'b11100101101101;     //325pi/512
  assign sin[326]  =  14'b11000101110100;     //326pi/512
  assign cos[326]  =  14'b11100101010110;     //326pi/512
  assign sin[327]  =  14'b11000101111111;     //327pi/512
  assign cos[327]  =  14'b11100100111111;     //327pi/512
  assign sin[328]  =  14'b11000110001001;     //328pi/512
  assign cos[328]  =  14'b11100100101001;     //328pi/512
  assign sin[329]  =  14'b11000110010100;     //329pi/512
  assign cos[329]  =  14'b11100100010010;     //329pi/512
  assign sin[330]  =  14'b11000110011111;     //330pi/512
  assign cos[330]  =  14'b11100011111011;     //330pi/512
  assign sin[331]  =  14'b11000110101010;     //331pi/512
  assign cos[331]  =  14'b11100011100101;     //331pi/512
  assign sin[332]  =  14'b11000110110101;     //332pi/512
  assign cos[332]  =  14'b11100011001110;     //332pi/512
  assign sin[333]  =  14'b11000111000001;     //333pi/512
  assign cos[333]  =  14'b11100010111000;     //333pi/512
  assign sin[334]  =  14'b11000111001100;     //334pi/512
  assign cos[334]  =  14'b11100010100010;     //334pi/512
  assign sin[335]  =  14'b11000111011000;     //335pi/512
  assign cos[335]  =  14'b11100010001011;     //335pi/512
  assign sin[336]  =  14'b11000111100100;     //336pi/512
  assign cos[336]  =  14'b11100001110101;     //336pi/512
  assign sin[337]  =  14'b11000111110000;     //337pi/512
  assign cos[337]  =  14'b11100001011111;     //337pi/512
  assign sin[338]  =  14'b11000111111100;     //338pi/512
  assign cos[338]  =  14'b11100001001001;     //338pi/512
  assign sin[339]  =  14'b11001000001000;     //339pi/512
  assign cos[339]  =  14'b11100000110011;     //339pi/512
  assign sin[340]  =  14'b11001000010100;     //340pi/512
  assign cos[340]  =  14'b11100000011101;     //340pi/512
  assign sin[341]  =  14'b11001000100001;     //341pi/512
  assign cos[341]  =  14'b11100000000111;     //341pi/512
  assign sin[342]  =  14'b11001000101101;     //342pi/512
  assign cos[342]  =  14'b11011111110010;     //342pi/512
  assign sin[343]  =  14'b11001000111010;     //343pi/512
  assign cos[343]  =  14'b11011111011100;     //343pi/512
  assign sin[344]  =  14'b11001001000111;     //344pi/512
  assign cos[344]  =  14'b11011111000110;     //344pi/512
  assign sin[345]  =  14'b11001001010100;     //345pi/512
  assign cos[345]  =  14'b11011110110001;     //345pi/512
  assign sin[346]  =  14'b11001001100001;     //346pi/512
  assign cos[346]  =  14'b11011110011011;     //346pi/512
  assign sin[347]  =  14'b11001001101110;     //347pi/512
  assign cos[347]  =  14'b11011110000110;     //347pi/512
  assign sin[348]  =  14'b11001001111011;     //348pi/512
  assign cos[348]  =  14'b11011101110001;     //348pi/512
  assign sin[349]  =  14'b11001010001001;     //349pi/512
  assign cos[349]  =  14'b11011101011011;     //349pi/512
  assign sin[350]  =  14'b11001010010111;     //350pi/512
  assign cos[350]  =  14'b11011101000110;     //350pi/512
  assign sin[351]  =  14'b11001010100100;     //351pi/512
  assign cos[351]  =  14'b11011100110001;     //351pi/512
  assign sin[352]  =  14'b11001010110010;     //352pi/512
  assign cos[352]  =  14'b11011100011100;     //352pi/512
  assign sin[353]  =  14'b11001011000000;     //353pi/512
  assign cos[353]  =  14'b11011100001000;     //353pi/512
  assign sin[354]  =  14'b11001011001110;     //354pi/512
  assign cos[354]  =  14'b11011011110011;     //354pi/512
  assign sin[355]  =  14'b11001011011101;     //355pi/512
  assign cos[355]  =  14'b11011011011110;     //355pi/512
  assign sin[356]  =  14'b11001011101011;     //356pi/512
  assign cos[356]  =  14'b11011011001001;     //356pi/512
  assign sin[357]  =  14'b11001011111010;     //357pi/512
  assign cos[357]  =  14'b11011010110101;     //357pi/512
  assign sin[358]  =  14'b11001100001000;     //358pi/512
  assign cos[358]  =  14'b11011010100001;     //358pi/512
  assign sin[359]  =  14'b11001100010111;     //359pi/512
  assign cos[359]  =  14'b11011010001100;     //359pi/512
  assign sin[360]  =  14'b11001100100110;     //360pi/512
  assign cos[360]  =  14'b11011001111000;     //360pi/512
  assign sin[361]  =  14'b11001100110101;     //361pi/512
  assign cos[361]  =  14'b11011001100100;     //361pi/512
  assign sin[362]  =  14'b11001101000100;     //362pi/512
  assign cos[362]  =  14'b11011001010000;     //362pi/512
  assign sin[363]  =  14'b11001101010100;     //363pi/512
  assign cos[363]  =  14'b11011000111100;     //363pi/512
  assign sin[364]  =  14'b11001101100011;     //364pi/512
  assign cos[364]  =  14'b11011000101000;     //364pi/512
  assign sin[365]  =  14'b11001101110010;     //365pi/512
  assign cos[365]  =  14'b11011000010100;     //365pi/512
  assign sin[366]  =  14'b11001110000010;     //366pi/512
  assign cos[366]  =  14'b11011000000001;     //366pi/512
  assign sin[367]  =  14'b11001110010010;     //367pi/512
  assign cos[367]  =  14'b11010111101101;     //367pi/512
  assign sin[368]  =  14'b11001110100010;     //368pi/512
  assign cos[368]  =  14'b11010111011010;     //368pi/512
  assign sin[369]  =  14'b11001110110010;     //369pi/512
  assign cos[369]  =  14'b11010111000110;     //369pi/512
  assign sin[370]  =  14'b11001111000010;     //370pi/512
  assign cos[370]  =  14'b11010110110011;     //370pi/512
  assign sin[371]  =  14'b11001111010010;     //371pi/512
  assign cos[371]  =  14'b11010110100000;     //371pi/512
  assign sin[372]  =  14'b11001111100010;     //372pi/512
  assign cos[372]  =  14'b11010110001101;     //372pi/512
  assign sin[373]  =  14'b11001111110011;     //373pi/512
  assign cos[373]  =  14'b11010101111010;     //373pi/512
  assign sin[374]  =  14'b11010000000100;     //374pi/512
  assign cos[374]  =  14'b11010101100111;     //374pi/512
  assign sin[375]  =  14'b11010000010100;     //375pi/512
  assign cos[375]  =  14'b11010101010100;     //375pi/512
  assign sin[376]  =  14'b11010000100101;     //376pi/512
  assign cos[376]  =  14'b11010101000001;     //376pi/512
  assign sin[377]  =  14'b11010000110110;     //377pi/512
  assign cos[377]  =  14'b11010100101111;     //377pi/512
  assign sin[378]  =  14'b11010001000111;     //378pi/512
  assign cos[378]  =  14'b11010100011100;     //378pi/512
  assign sin[379]  =  14'b11010001011000;     //379pi/512
  assign cos[379]  =  14'b11010100001010;     //379pi/512
  assign sin[380]  =  14'b11010001101001;     //380pi/512
  assign cos[380]  =  14'b11010011111000;     //380pi/512
  assign sin[381]  =  14'b11010001111011;     //381pi/512
  assign cos[381]  =  14'b11010011100101;     //381pi/512
  assign sin[382]  =  14'b11010010001100;     //382pi/512
  assign cos[382]  =  14'b11010011010011;     //382pi/512
  assign sin[383]  =  14'b11010010011110;     //383pi/512
  assign cos[383]  =  14'b11010011000010;     //383pi/512
  assign sin[384]  =  14'b11010010110000;     //384pi/512
  assign cos[384]  =  14'b11010010110000;     //384pi/512
  assign sin[385]  =  14'b11010011000010;     //385pi/512
  assign cos[385]  =  14'b11010010011110;     //385pi/512
  assign sin[386]  =  14'b11010011010011;     //386pi/512
  assign cos[386]  =  14'b11010010001100;     //386pi/512
  assign sin[387]  =  14'b11010011100101;     //387pi/512
  assign cos[387]  =  14'b11010001111011;     //387pi/512
  assign sin[388]  =  14'b11010011111000;     //388pi/512
  assign cos[388]  =  14'b11010001101001;     //388pi/512
  assign sin[389]  =  14'b11010100001010;     //389pi/512
  assign cos[389]  =  14'b11010001011000;     //389pi/512
  assign sin[390]  =  14'b11010100011100;     //390pi/512
  assign cos[390]  =  14'b11010001000111;     //390pi/512
  assign sin[391]  =  14'b11010100101111;     //391pi/512
  assign cos[391]  =  14'b11010000110110;     //391pi/512
  assign sin[392]  =  14'b11010101000001;     //392pi/512
  assign cos[392]  =  14'b11010000100101;     //392pi/512
  assign sin[393]  =  14'b11010101010100;     //393pi/512
  assign cos[393]  =  14'b11010000010100;     //393pi/512
  assign sin[394]  =  14'b11010101100111;     //394pi/512
  assign cos[394]  =  14'b11010000000100;     //394pi/512
  assign sin[395]  =  14'b11010101111010;     //395pi/512
  assign cos[395]  =  14'b11001111110011;     //395pi/512
  assign sin[396]  =  14'b11010110001101;     //396pi/512
  assign cos[396]  =  14'b11001111100010;     //396pi/512
  assign sin[397]  =  14'b11010110100000;     //397pi/512
  assign cos[397]  =  14'b11001111010010;     //397pi/512
  assign sin[398]  =  14'b11010110110011;     //398pi/512
  assign cos[398]  =  14'b11001111000010;     //398pi/512
  assign sin[399]  =  14'b11010111000110;     //399pi/512
  assign cos[399]  =  14'b11001110110010;     //399pi/512
  assign sin[400]  =  14'b11010111011010;     //400pi/512
  assign cos[400]  =  14'b11001110100010;     //400pi/512
  assign sin[401]  =  14'b11010111101101;     //401pi/512
  assign cos[401]  =  14'b11001110010010;     //401pi/512
  assign sin[402]  =  14'b11011000000001;     //402pi/512
  assign cos[402]  =  14'b11001110000010;     //402pi/512
  assign sin[403]  =  14'b11011000010100;     //403pi/512
  assign cos[403]  =  14'b11001101110010;     //403pi/512
  assign sin[404]  =  14'b11011000101000;     //404pi/512
  assign cos[404]  =  14'b11001101100011;     //404pi/512
  assign sin[405]  =  14'b11011000111100;     //405pi/512
  assign cos[405]  =  14'b11001101010100;     //405pi/512
  assign sin[406]  =  14'b11011001010000;     //406pi/512
  assign cos[406]  =  14'b11001101000100;     //406pi/512
  assign sin[407]  =  14'b11011001100100;     //407pi/512
  assign cos[407]  =  14'b11001100110101;     //407pi/512
  assign sin[408]  =  14'b11011001111000;     //408pi/512
  assign cos[408]  =  14'b11001100100110;     //408pi/512
  assign sin[409]  =  14'b11011010001100;     //409pi/512
  assign cos[409]  =  14'b11001100010111;     //409pi/512
  assign sin[410]  =  14'b11011010100001;     //410pi/512
  assign cos[410]  =  14'b11001100001000;     //410pi/512
  assign sin[411]  =  14'b11011010110101;     //411pi/512
  assign cos[411]  =  14'b11001011111010;     //411pi/512
  assign sin[412]  =  14'b11011011001001;     //412pi/512
  assign cos[412]  =  14'b11001011101011;     //412pi/512
  assign sin[413]  =  14'b11011011011110;     //413pi/512
  assign cos[413]  =  14'b11001011011101;     //413pi/512
  assign sin[414]  =  14'b11011011110011;     //414pi/512
  assign cos[414]  =  14'b11001011001110;     //414pi/512
  assign sin[415]  =  14'b11011100001000;     //415pi/512
  assign cos[415]  =  14'b11001011000000;     //415pi/512
  assign sin[416]  =  14'b11011100011100;     //416pi/512
  assign cos[416]  =  14'b11001010110010;     //416pi/512
  assign sin[417]  =  14'b11011100110001;     //417pi/512
  assign cos[417]  =  14'b11001010100100;     //417pi/512
  assign sin[418]  =  14'b11011101000110;     //418pi/512
  assign cos[418]  =  14'b11001010010111;     //418pi/512
  assign sin[419]  =  14'b11011101011011;     //419pi/512
  assign cos[419]  =  14'b11001010001001;     //419pi/512
  assign sin[420]  =  14'b11011101110001;     //420pi/512
  assign cos[420]  =  14'b11001001111011;     //420pi/512
  assign sin[421]  =  14'b11011110000110;     //421pi/512
  assign cos[421]  =  14'b11001001101110;     //421pi/512
  assign sin[422]  =  14'b11011110011011;     //422pi/512
  assign cos[422]  =  14'b11001001100001;     //422pi/512
  assign sin[423]  =  14'b11011110110001;     //423pi/512
  assign cos[423]  =  14'b11001001010100;     //423pi/512
  assign sin[424]  =  14'b11011111000110;     //424pi/512
  assign cos[424]  =  14'b11001001000111;     //424pi/512
  assign sin[425]  =  14'b11011111011100;     //425pi/512
  assign cos[425]  =  14'b11001000111010;     //425pi/512
  assign sin[426]  =  14'b11011111110010;     //426pi/512
  assign cos[426]  =  14'b11001000101101;     //426pi/512
  assign sin[427]  =  14'b11100000000111;     //427pi/512
  assign cos[427]  =  14'b11001000100001;     //427pi/512
  assign sin[428]  =  14'b11100000011101;     //428pi/512
  assign cos[428]  =  14'b11001000010100;     //428pi/512
  assign sin[429]  =  14'b11100000110011;     //429pi/512
  assign cos[429]  =  14'b11001000001000;     //429pi/512
  assign sin[430]  =  14'b11100001001001;     //430pi/512
  assign cos[430]  =  14'b11000111111100;     //430pi/512
  assign sin[431]  =  14'b11100001011111;     //431pi/512
  assign cos[431]  =  14'b11000111110000;     //431pi/512
  assign sin[432]  =  14'b11100001110101;     //432pi/512
  assign cos[432]  =  14'b11000111100100;     //432pi/512
  assign sin[433]  =  14'b11100010001011;     //433pi/512
  assign cos[433]  =  14'b11000111011000;     //433pi/512
  assign sin[434]  =  14'b11100010100010;     //434pi/512
  assign cos[434]  =  14'b11000111001100;     //434pi/512
  assign sin[435]  =  14'b11100010111000;     //435pi/512
  assign cos[435]  =  14'b11000111000001;     //435pi/512
  assign sin[436]  =  14'b11100011001110;     //436pi/512
  assign cos[436]  =  14'b11000110110101;     //436pi/512
  assign sin[437]  =  14'b11100011100101;     //437pi/512
  assign cos[437]  =  14'b11000110101010;     //437pi/512
  assign sin[438]  =  14'b11100011111011;     //438pi/512
  assign cos[438]  =  14'b11000110011111;     //438pi/512
  assign sin[439]  =  14'b11100100010010;     //439pi/512
  assign cos[439]  =  14'b11000110010100;     //439pi/512
  assign sin[440]  =  14'b11100100101001;     //440pi/512
  assign cos[440]  =  14'b11000110001001;     //440pi/512
  assign sin[441]  =  14'b11100100111111;     //441pi/512
  assign cos[441]  =  14'b11000101111111;     //441pi/512
  assign sin[442]  =  14'b11100101010110;     //442pi/512
  assign cos[442]  =  14'b11000101110100;     //442pi/512
  assign sin[443]  =  14'b11100101101101;     //443pi/512
  assign cos[443]  =  14'b11000101101010;     //443pi/512
  assign sin[444]  =  14'b11100110000100;     //444pi/512
  assign cos[444]  =  14'b11000101011111;     //444pi/512
  assign sin[445]  =  14'b11100110011011;     //445pi/512
  assign cos[445]  =  14'b11000101010101;     //445pi/512
  assign sin[446]  =  14'b11100110110010;     //446pi/512
  assign cos[446]  =  14'b11000101001011;     //446pi/512
  assign sin[447]  =  14'b11100111001001;     //447pi/512
  assign cos[447]  =  14'b11000101000001;     //447pi/512
  assign sin[448]  =  14'b11100111100001;     //448pi/512
  assign cos[448]  =  14'b11000100111000;     //448pi/512
  assign sin[449]  =  14'b11100111111000;     //449pi/512
  assign cos[449]  =  14'b11000100101110;     //449pi/512
  assign sin[450]  =  14'b11101000001111;     //450pi/512
  assign cos[450]  =  14'b11000100100101;     //450pi/512
  assign sin[451]  =  14'b11101000100110;     //451pi/512
  assign cos[451]  =  14'b11000100011100;     //451pi/512
  assign sin[452]  =  14'b11101000111110;     //452pi/512
  assign cos[452]  =  14'b11000100010010;     //452pi/512
  assign sin[453]  =  14'b11101001010101;     //453pi/512
  assign cos[453]  =  14'b11000100001001;     //453pi/512
  assign sin[454]  =  14'b11101001101101;     //454pi/512
  assign cos[454]  =  14'b11000100000001;     //454pi/512
  assign sin[455]  =  14'b11101010000100;     //455pi/512
  assign cos[455]  =  14'b11000011111000;     //455pi/512
  assign sin[456]  =  14'b11101010011100;     //456pi/512
  assign cos[456]  =  14'b11000011101111;     //456pi/512
  assign sin[457]  =  14'b11101010110100;     //457pi/512
  assign cos[457]  =  14'b11000011100111;     //457pi/512
  assign sin[458]  =  14'b11101011001100;     //458pi/512
  assign cos[458]  =  14'b11000011011111;     //458pi/512
  assign sin[459]  =  14'b11101011100011;     //459pi/512
  assign cos[459]  =  14'b11000011010111;     //459pi/512
  assign sin[460]  =  14'b11101011111011;     //460pi/512
  assign cos[460]  =  14'b11000011001111;     //460pi/512
  assign sin[461]  =  14'b11101100010011;     //461pi/512
  assign cos[461]  =  14'b11000011000111;     //461pi/512
  assign sin[462]  =  14'b11101100101011;     //462pi/512
  assign cos[462]  =  14'b11000010111111;     //462pi/512
  assign sin[463]  =  14'b11101101000011;     //463pi/512
  assign cos[463]  =  14'b11000010111000;     //463pi/512
  assign sin[464]  =  14'b11101101011011;     //464pi/512
  assign cos[464]  =  14'b11000010110000;     //464pi/512
  assign sin[465]  =  14'b11101101110011;     //465pi/512
  assign cos[465]  =  14'b11000010101001;     //465pi/512
  assign sin[466]  =  14'b11101110001011;     //466pi/512
  assign cos[466]  =  14'b11000010100010;     //466pi/512
  assign sin[467]  =  14'b11101110100011;     //467pi/512
  assign cos[467]  =  14'b11000010011011;     //467pi/512
  assign sin[468]  =  14'b11101110111100;     //468pi/512
  assign cos[468]  =  14'b11000010010100;     //468pi/512
  assign sin[469]  =  14'b11101111010100;     //469pi/512
  assign cos[469]  =  14'b11000010001110;     //469pi/512
  assign sin[470]  =  14'b11101111101100;     //470pi/512
  assign cos[470]  =  14'b11000010000111;     //470pi/512
  assign sin[471]  =  14'b11110000000100;     //471pi/512
  assign cos[471]  =  14'b11000010000001;     //471pi/512
  assign sin[472]  =  14'b11110000011101;     //472pi/512
  assign cos[472]  =  14'b11000001111011;     //472pi/512
  assign sin[473]  =  14'b11110000110101;     //473pi/512
  assign cos[473]  =  14'b11000001110101;     //473pi/512
  assign sin[474]  =  14'b11110001001110;     //474pi/512
  assign cos[474]  =  14'b11000001101111;     //474pi/512
  assign sin[475]  =  14'b11110001100110;     //475pi/512
  assign cos[475]  =  14'b11000001101001;     //475pi/512
  assign sin[476]  =  14'b11110001111111;     //476pi/512
  assign cos[476]  =  14'b11000001100100;     //476pi/512
  assign sin[477]  =  14'b11110010010111;     //477pi/512
  assign cos[477]  =  14'b11000001011110;     //477pi/512
  assign sin[478]  =  14'b11110010110000;     //478pi/512
  assign cos[478]  =  14'b11000001011001;     //478pi/512
  assign sin[479]  =  14'b11110011001000;     //479pi/512
  assign cos[479]  =  14'b11000001010100;     //479pi/512
  assign sin[480]  =  14'b11110011100001;     //480pi/512
  assign cos[480]  =  14'b11000001001111;     //480pi/512
  assign sin[481]  =  14'b11110011111010;     //481pi/512
  assign cos[481]  =  14'b11000001001010;     //481pi/512
  assign sin[482]  =  14'b11110100010010;     //482pi/512
  assign cos[482]  =  14'b11000001000101;     //482pi/512
  assign sin[483]  =  14'b11110100101011;     //483pi/512
  assign cos[483]  =  14'b11000001000001;     //483pi/512
  assign sin[484]  =  14'b11110101000100;     //484pi/512
  assign cos[484]  =  14'b11000000111100;     //484pi/512
  assign sin[485]  =  14'b11110101011101;     //485pi/512
  assign cos[485]  =  14'b11000000111000;     //485pi/512
  assign sin[486]  =  14'b11110101110101;     //486pi/512
  assign cos[486]  =  14'b11000000110100;     //486pi/512
  assign sin[487]  =  14'b11110110001110;     //487pi/512
  assign cos[487]  =  14'b11000000110000;     //487pi/512
  assign sin[488]  =  14'b11110110100111;     //488pi/512
  assign cos[488]  =  14'b11000000101100;     //488pi/512
  assign sin[489]  =  14'b11110111000000;     //489pi/512
  assign cos[489]  =  14'b11000000101001;     //489pi/512
  assign sin[490]  =  14'b11110111011001;     //490pi/512
  assign cos[490]  =  14'b11000000100101;     //490pi/512
  assign sin[491]  =  14'b11110111110010;     //491pi/512
  assign cos[491]  =  14'b11000000100010;     //491pi/512
  assign sin[492]  =  14'b11111000001011;     //492pi/512
  assign cos[492]  =  14'b11000000011111;     //492pi/512
  assign sin[493]  =  14'b11111000100100;     //493pi/512
  assign cos[493]  =  14'b11000000011100;     //493pi/512
  assign sin[494]  =  14'b11111000111101;     //494pi/512
  assign cos[494]  =  14'b11000000011001;     //494pi/512
  assign sin[495]  =  14'b11111001010110;     //495pi/512
  assign cos[495]  =  14'b11000000010110;     //495pi/512
  assign sin[496]  =  14'b11111001101111;     //496pi/512
  assign cos[496]  =  14'b11000000010100;     //496pi/512
  assign sin[497]  =  14'b11111010001000;     //497pi/512
  assign cos[497]  =  14'b11000000010001;     //497pi/512
  assign sin[498]  =  14'b11111010100001;     //498pi/512
  assign cos[498]  =  14'b11000000001111;     //498pi/512
  assign sin[499]  =  14'b11111010111010;     //499pi/512
  assign cos[499]  =  14'b11000000001101;     //499pi/512
  assign sin[500]  =  14'b11111011010011;     //500pi/512
  assign cos[500]  =  14'b11000000001011;     //500pi/512
  assign sin[501]  =  14'b11111011101100;     //501pi/512
  assign cos[501]  =  14'b11000000001001;     //501pi/512
  assign sin[502]  =  14'b11111100000101;     //502pi/512
  assign cos[502]  =  14'b11000000001000;     //502pi/512
  assign sin[503]  =  14'b11111100011110;     //503pi/512
  assign cos[503]  =  14'b11000000000110;     //503pi/512
  assign sin[504]  =  14'b11111100110111;     //504pi/512
  assign cos[504]  =  14'b11000000000101;     //504pi/512
  assign sin[505]  =  14'b11111101010000;     //505pi/512
  assign cos[505]  =  14'b11000000000100;     //505pi/512
  assign sin[506]  =  14'b11111101101001;     //506pi/512
  assign cos[506]  =  14'b11000000000011;     //506pi/512
  assign sin[507]  =  14'b11111110000010;     //507pi/512
  assign cos[507]  =  14'b11000000000010;     //507pi/512
  assign sin[508]  =  14'b11111110011011;     //508pi/512
  assign cos[508]  =  14'b11000000000001;     //508pi/512
  assign sin[509]  =  14'b11111110110101;     //509pi/512
  assign cos[509]  =  14'b11000000000001;     //509pi/512
  assign sin[510]  =  14'b11111111001110;     //510pi/512
  assign cos[510]  =  14'b11000000000000;     //510pi/512
  assign sin[511]  =  14'b11111111100111;     //511pi/512
  assign cos[511]  =  14'b11000000000000;     //511pi/512

  assign sin2[0]  =  14'b00000000000000;     //0pi/512
  assign cos2[0]  =  14'b01000000000000;     //0pi/512
  assign sin2[1]  =  14'b11111111101100;     //1pi/512
  assign cos2[1]  =  14'b00111111111111;     //1pi/512
  assign sin2[2]  =  14'b11111111011000;     //2pi/512
  assign cos2[2]  =  14'b00111111111111;     //2pi/512
  assign sin2[3]  =  14'b11111111000100;     //3pi/512
  assign cos2[3]  =  14'b00111111111111;     //3pi/512
  assign sin2[4]  =  14'b11111110110000;     //4pi/512
  assign cos2[4]  =  14'b00111111111111;     //4pi/512
  assign sin2[5]  =  14'b11111110011011;     //5pi/512
  assign cos2[5]  =  14'b00111111111110;     //5pi/512
  assign sin2[6]  =  14'b11111110000111;     //6pi/512
  assign cos2[6]  =  14'b00111111111110;     //6pi/512
  assign sin2[7]  =  14'b11111101110011;     //7pi/512
  assign cos2[7]  =  14'b00111111111101;     //7pi/512
  assign sin2[8]  =  14'b11111101011111;     //8pi/512
  assign cos2[8]  =  14'b00111111111100;     //8pi/512
  assign sin2[9]  =  14'b11111101001011;     //9pi/512
  assign cos2[9]  =  14'b00111111111100;     //9pi/512
  assign sin2[10]  =  14'b11111100110111;     //10pi/512
  assign cos2[10]  =  14'b00111111111011;     //10pi/512
  assign sin2[11]  =  14'b11111100100011;     //11pi/512
  assign cos2[11]  =  14'b00111111111010;     //11pi/512
  assign sin2[12]  =  14'b11111100001111;     //12pi/512
  assign cos2[12]  =  14'b00111111111000;     //12pi/512
  assign sin2[13]  =  14'b11111011111011;     //13pi/512
  assign cos2[13]  =  14'b00111111110111;     //13pi/512
  assign sin2[14]  =  14'b11111011100111;     //14pi/512
  assign cos2[14]  =  14'b00111111110110;     //14pi/512
  assign sin2[15]  =  14'b11111011010011;     //15pi/512
  assign cos2[15]  =  14'b00111111110100;     //15pi/512
  assign sin2[16]  =  14'b11111010111111;     //16pi/512
  assign cos2[16]  =  14'b00111111110011;     //16pi/512
  assign sin2[17]  =  14'b11111010101011;     //17pi/512
  assign cos2[17]  =  14'b00111111110001;     //17pi/512
  assign sin2[18]  =  14'b11111010010111;     //18pi/512
  assign cos2[18]  =  14'b00111111110000;     //18pi/512
  assign sin2[19]  =  14'b11111010000011;     //19pi/512
  assign cos2[19]  =  14'b00111111101110;     //19pi/512
  assign sin2[20]  =  14'b11111001101111;     //20pi/512
  assign cos2[20]  =  14'b00111111101100;     //20pi/512
  assign sin2[21]  =  14'b11111001011011;     //21pi/512
  assign cos2[21]  =  14'b00111111101010;     //21pi/512
  assign sin2[22]  =  14'b11111001000111;     //22pi/512
  assign cos2[22]  =  14'b00111111101000;     //22pi/512
  assign sin2[23]  =  14'b11111000110011;     //23pi/512
  assign cos2[23]  =  14'b00111111100101;     //23pi/512
  assign sin2[24]  =  14'b11111000011111;     //24pi/512
  assign cos2[24]  =  14'b00111111100011;     //24pi/512
  assign sin2[25]  =  14'b11111000001011;     //25pi/512
  assign cos2[25]  =  14'b00111111100001;     //25pi/512
  assign sin2[26]  =  14'b11110111110111;     //26pi/512
  assign cos2[26]  =  14'b00111111011110;     //26pi/512
  assign sin2[27]  =  14'b11110111100011;     //27pi/512
  assign cos2[27]  =  14'b00111111011100;     //27pi/512
  assign sin2[28]  =  14'b11110111001111;     //28pi/512
  assign cos2[28]  =  14'b00111111011001;     //28pi/512
  assign sin2[29]  =  14'b11110110111011;     //29pi/512
  assign cos2[29]  =  14'b00111111010110;     //29pi/512
  assign sin2[30]  =  14'b11110110100111;     //30pi/512
  assign cos2[30]  =  14'b00111111010011;     //30pi/512
  assign sin2[31]  =  14'b11110110010011;     //31pi/512
  assign cos2[31]  =  14'b00111111010000;     //31pi/512
  assign sin2[32]  =  14'b11110101111111;     //32pi/512
  assign cos2[32]  =  14'b00111111001101;     //32pi/512
  assign sin2[33]  =  14'b11110101101011;     //33pi/512
  assign cos2[33]  =  14'b00111111001010;     //33pi/512
  assign sin2[34]  =  14'b11110101011000;     //34pi/512
  assign cos2[34]  =  14'b00111111000111;     //34pi/512
  assign sin2[35]  =  14'b11110101000100;     //35pi/512
  assign cos2[35]  =  14'b00111111000011;     //35pi/512
  assign sin2[36]  =  14'b11110100110000;     //36pi/512
  assign cos2[36]  =  14'b00111111000000;     //36pi/512
  assign sin2[37]  =  14'b11110100011100;     //37pi/512
  assign cos2[37]  =  14'b00111110111100;     //37pi/512
  assign sin2[38]  =  14'b11110100001000;     //38pi/512
  assign cos2[38]  =  14'b00111110111000;     //38pi/512
  assign sin2[39]  =  14'b11110011110101;     //39pi/512
  assign cos2[39]  =  14'b00111110110101;     //39pi/512
  assign sin2[40]  =  14'b11110011100001;     //40pi/512
  assign cos2[40]  =  14'b00111110110001;     //40pi/512
  assign sin2[41]  =  14'b11110011001101;     //41pi/512
  assign cos2[41]  =  14'b00111110101101;     //41pi/512
  assign sin2[42]  =  14'b11110010111010;     //42pi/512
  assign cos2[42]  =  14'b00111110101001;     //42pi/512
  assign sin2[43]  =  14'b11110010100110;     //43pi/512
  assign cos2[43]  =  14'b00111110100101;     //43pi/512
  assign sin2[44]  =  14'b11110010010010;     //44pi/512
  assign cos2[44]  =  14'b00111110100000;     //44pi/512
  assign sin2[45]  =  14'b11110001111111;     //45pi/512
  assign cos2[45]  =  14'b00111110011100;     //45pi/512
  assign sin2[46]  =  14'b11110001101011;     //46pi/512
  assign cos2[46]  =  14'b00111110011000;     //46pi/512
  assign sin2[47]  =  14'b11110001010111;     //47pi/512
  assign cos2[47]  =  14'b00111110010011;     //47pi/512
  assign sin2[48]  =  14'b11110001000100;     //48pi/512
  assign cos2[48]  =  14'b00111110001110;     //48pi/512
  assign sin2[49]  =  14'b11110000110000;     //49pi/512
  assign cos2[49]  =  14'b00111110001010;     //49pi/512
  assign sin2[50]  =  14'b11110000011101;     //50pi/512
  assign cos2[50]  =  14'b00111110000101;     //50pi/512
  assign sin2[51]  =  14'b11110000001001;     //51pi/512
  assign cos2[51]  =  14'b00111110000000;     //51pi/512
  assign sin2[52]  =  14'b11101111110110;     //52pi/512
  assign cos2[52]  =  14'b00111101111011;     //52pi/512
  assign sin2[53]  =  14'b11101111100010;     //53pi/512
  assign cos2[53]  =  14'b00111101110110;     //53pi/512
  assign sin2[54]  =  14'b11101111001111;     //54pi/512
  assign cos2[54]  =  14'b00111101110000;     //54pi/512
  assign sin2[55]  =  14'b11101110111100;     //55pi/512
  assign cos2[55]  =  14'b00111101101011;     //55pi/512
  assign sin2[56]  =  14'b11101110101000;     //56pi/512
  assign cos2[56]  =  14'b00111101100110;     //56pi/512
  assign sin2[57]  =  14'b11101110010101;     //57pi/512
  assign cos2[57]  =  14'b00111101100000;     //57pi/512
  assign sin2[58]  =  14'b11101110000010;     //58pi/512
  assign cos2[58]  =  14'b00111101011011;     //58pi/512
  assign sin2[59]  =  14'b11101101101110;     //59pi/512
  assign cos2[59]  =  14'b00111101010101;     //59pi/512
  assign sin2[60]  =  14'b11101101011011;     //60pi/512
  assign cos2[60]  =  14'b00111101001111;     //60pi/512
  assign sin2[61]  =  14'b11101101001000;     //61pi/512
  assign cos2[61]  =  14'b00111101001001;     //61pi/512
  assign sin2[62]  =  14'b11101100110101;     //62pi/512
  assign cos2[62]  =  14'b00111101000011;     //62pi/512
  assign sin2[63]  =  14'b11101100100001;     //63pi/512
  assign cos2[63]  =  14'b00111100111101;     //63pi/512
  assign sin2[64]  =  14'b11101100001110;     //64pi/512
  assign cos2[64]  =  14'b00111100110111;     //64pi/512
  assign sin2[65]  =  14'b11101011111011;     //65pi/512
  assign cos2[65]  =  14'b00111100110001;     //65pi/512
  assign sin2[66]  =  14'b11101011101000;     //66pi/512
  assign cos2[66]  =  14'b00111100101010;     //66pi/512
  assign sin2[67]  =  14'b11101011010101;     //67pi/512
  assign cos2[67]  =  14'b00111100100100;     //67pi/512
  assign sin2[68]  =  14'b11101011000010;     //68pi/512
  assign cos2[68]  =  14'b00111100011101;     //68pi/512
  assign sin2[69]  =  14'b11101010101111;     //69pi/512
  assign cos2[69]  =  14'b00111100010111;     //69pi/512
  assign sin2[70]  =  14'b11101010011100;     //70pi/512
  assign cos2[70]  =  14'b00111100010000;     //70pi/512
  assign sin2[71]  =  14'b11101010001001;     //71pi/512
  assign cos2[71]  =  14'b00111100001001;     //71pi/512
  assign sin2[72]  =  14'b11101001110110;     //72pi/512
  assign cos2[72]  =  14'b00111100000010;     //72pi/512
  assign sin2[73]  =  14'b11101001100011;     //73pi/512
  assign cos2[73]  =  14'b00111011111011;     //73pi/512
  assign sin2[74]  =  14'b11101001010001;     //74pi/512
  assign cos2[74]  =  14'b00111011110100;     //74pi/512
  assign sin2[75]  =  14'b11101000111110;     //75pi/512
  assign cos2[75]  =  14'b00111011101101;     //75pi/512
  assign sin2[76]  =  14'b11101000101011;     //76pi/512
  assign cos2[76]  =  14'b00111011100110;     //76pi/512
  assign sin2[77]  =  14'b11101000011000;     //77pi/512
  assign cos2[77]  =  14'b00111011011110;     //77pi/512
  assign sin2[78]  =  14'b11101000000110;     //78pi/512
  assign cos2[78]  =  14'b00111011010111;     //78pi/512
  assign sin2[79]  =  14'b11100111110011;     //79pi/512
  assign cos2[79]  =  14'b00111011001111;     //79pi/512
  assign sin2[80]  =  14'b11100111100001;     //80pi/512
  assign cos2[80]  =  14'b00111011001000;     //80pi/512
  assign sin2[81]  =  14'b11100111001110;     //81pi/512
  assign cos2[81]  =  14'b00111011000000;     //81pi/512
  assign sin2[82]  =  14'b11100110111011;     //82pi/512
  assign cos2[82]  =  14'b00111010111000;     //82pi/512
  assign sin2[83]  =  14'b11100110101001;     //83pi/512
  assign cos2[83]  =  14'b00111010110000;     //83pi/512
  assign sin2[84]  =  14'b11100110010111;     //84pi/512
  assign cos2[84]  =  14'b00111010101000;     //84pi/512
  assign sin2[85]  =  14'b11100110000100;     //85pi/512
  assign cos2[85]  =  14'b00111010100000;     //85pi/512
  assign sin2[86]  =  14'b11100101110010;     //86pi/512
  assign cos2[86]  =  14'b00111010011000;     //86pi/512
  assign sin2[87]  =  14'b11100101011111;     //87pi/512
  assign cos2[87]  =  14'b00111010010000;     //87pi/512
  assign sin2[88]  =  14'b11100101001101;     //88pi/512
  assign cos2[88]  =  14'b00111010000111;     //88pi/512
  assign sin2[89]  =  14'b11100100111011;     //89pi/512
  assign cos2[89]  =  14'b00111001111111;     //89pi/512
  assign sin2[90]  =  14'b11100100101001;     //90pi/512
  assign cos2[90]  =  14'b00111001110110;     //90pi/512
  assign sin2[91]  =  14'b11100100010111;     //91pi/512
  assign cos2[91]  =  14'b00111001101110;     //91pi/512
  assign sin2[92]  =  14'b11100100000100;     //92pi/512
  assign cos2[92]  =  14'b00111001100101;     //92pi/512
  assign sin2[93]  =  14'b11100011110010;     //93pi/512
  assign cos2[93]  =  14'b00111001011100;     //93pi/512
  assign sin2[94]  =  14'b11100011100000;     //94pi/512
  assign cos2[94]  =  14'b00111001010011;     //94pi/512
  assign sin2[95]  =  14'b11100011001110;     //95pi/512
  assign cos2[95]  =  14'b00111001001010;     //95pi/512
  assign sin2[96]  =  14'b11100010111100;     //96pi/512
  assign cos2[96]  =  14'b00111001000001;     //96pi/512
  assign sin2[97]  =  14'b11100010101011;     //97pi/512
  assign cos2[97]  =  14'b00111000111000;     //97pi/512
  assign sin2[98]  =  14'b11100010011001;     //98pi/512
  assign cos2[98]  =  14'b00111000101111;     //98pi/512
  assign sin2[99]  =  14'b11100010000111;     //99pi/512
  assign cos2[99]  =  14'b00111000100101;     //99pi/512
  assign sin2[100]  =  14'b11100001110101;     //100pi/512
  assign cos2[100]  =  14'b00111000011100;     //100pi/512
  assign sin2[101]  =  14'b11100001100011;     //101pi/512
  assign cos2[101]  =  14'b00111000010010;     //101pi/512
  assign sin2[102]  =  14'b11100001010010;     //102pi/512
  assign cos2[102]  =  14'b00111000001001;     //102pi/512
  assign sin2[103]  =  14'b11100001000000;     //103pi/512
  assign cos2[103]  =  14'b00110111111111;     //103pi/512
  assign sin2[104]  =  14'b11100000101111;     //104pi/512
  assign cos2[104]  =  14'b00110111110101;     //104pi/512
  assign sin2[105]  =  14'b11100000011101;     //105pi/512
  assign cos2[105]  =  14'b00110111101011;     //105pi/512
  assign sin2[106]  =  14'b11100000001100;     //106pi/512
  assign cos2[106]  =  14'b00110111100001;     //106pi/512
  assign sin2[107]  =  14'b11011111111010;     //107pi/512
  assign cos2[107]  =  14'b00110111010111;     //107pi/512
  assign sin2[108]  =  14'b11011111101001;     //108pi/512
  assign cos2[108]  =  14'b00110111001101;     //108pi/512
  assign sin2[109]  =  14'b11011111011000;     //109pi/512
  assign cos2[109]  =  14'b00110111000011;     //109pi/512
  assign sin2[110]  =  14'b11011111000110;     //110pi/512
  assign cos2[110]  =  14'b00110110111001;     //110pi/512
  assign sin2[111]  =  14'b11011110110101;     //111pi/512
  assign cos2[111]  =  14'b00110110101110;     //111pi/512
  assign sin2[112]  =  14'b11011110100100;     //112pi/512
  assign cos2[112]  =  14'b00110110100100;     //112pi/512
  assign sin2[113]  =  14'b11011110010011;     //113pi/512
  assign cos2[113]  =  14'b00110110011001;     //113pi/512
  assign sin2[114]  =  14'b11011110000010;     //114pi/512
  assign cos2[114]  =  14'b00110110001111;     //114pi/512
  assign sin2[115]  =  14'b11011101110001;     //115pi/512
  assign cos2[115]  =  14'b00110110000100;     //115pi/512
  assign sin2[116]  =  14'b11011101100000;     //116pi/512
  assign cos2[116]  =  14'b00110101111001;     //116pi/512
  assign sin2[117]  =  14'b11011101001111;     //117pi/512
  assign cos2[117]  =  14'b00110101101110;     //117pi/512
  assign sin2[118]  =  14'b11011100111110;     //118pi/512
  assign cos2[118]  =  14'b00110101100011;     //118pi/512
  assign sin2[119]  =  14'b11011100101101;     //119pi/512
  assign cos2[119]  =  14'b00110101011000;     //119pi/512
  assign sin2[120]  =  14'b11011100011100;     //120pi/512
  assign cos2[120]  =  14'b00110101001101;     //120pi/512
  assign sin2[121]  =  14'b11011100001100;     //121pi/512
  assign cos2[121]  =  14'b00110101000010;     //121pi/512
  assign sin2[122]  =  14'b11011011111011;     //122pi/512
  assign cos2[122]  =  14'b00110100110111;     //122pi/512
  assign sin2[123]  =  14'b11011011101010;     //123pi/512
  assign cos2[123]  =  14'b00110100101011;     //123pi/512
  assign sin2[124]  =  14'b11011011011010;     //124pi/512
  assign cos2[124]  =  14'b00110100100000;     //124pi/512
  assign sin2[125]  =  14'b11011011001001;     //125pi/512
  assign cos2[125]  =  14'b00110100010100;     //125pi/512
  assign sin2[126]  =  14'b11011010111001;     //126pi/512
  assign cos2[126]  =  14'b00110100001001;     //126pi/512
  assign sin2[127]  =  14'b11011010101001;     //127pi/512
  assign cos2[127]  =  14'b00110011111101;     //127pi/512
  assign sin2[128]  =  14'b11011010011000;     //128pi/512
  assign cos2[128]  =  14'b00110011110001;     //128pi/512
  assign sin2[129]  =  14'b11011010001000;     //129pi/512
  assign cos2[129]  =  14'b00110011100101;     //129pi/512
  assign sin2[130]  =  14'b11011001111000;     //130pi/512
  assign cos2[130]  =  14'b00110011011001;     //130pi/512
  assign sin2[131]  =  14'b11011001101000;     //131pi/512
  assign cos2[131]  =  14'b00110011001101;     //131pi/512
  assign sin2[132]  =  14'b11011001011000;     //132pi/512
  assign cos2[132]  =  14'b00110011000001;     //132pi/512
  assign sin2[133]  =  14'b11011001001000;     //133pi/512
  assign cos2[133]  =  14'b00110010110101;     //133pi/512
  assign sin2[134]  =  14'b11011000111000;     //134pi/512
  assign cos2[134]  =  14'b00110010101001;     //134pi/512
  assign sin2[135]  =  14'b11011000101000;     //135pi/512
  assign cos2[135]  =  14'b00110010011101;     //135pi/512
  assign sin2[136]  =  14'b11011000011000;     //136pi/512
  assign cos2[136]  =  14'b00110010010000;     //136pi/512
  assign sin2[137]  =  14'b11011000001000;     //137pi/512
  assign cos2[137]  =  14'b00110010000100;     //137pi/512
  assign sin2[138]  =  14'b11010111111001;     //138pi/512
  assign cos2[138]  =  14'b00110001110111;     //138pi/512
  assign sin2[139]  =  14'b11010111101001;     //139pi/512
  assign cos2[139]  =  14'b00110001101010;     //139pi/512
  assign sin2[140]  =  14'b11010111011010;     //140pi/512
  assign cos2[140]  =  14'b00110001011110;     //140pi/512
  assign sin2[141]  =  14'b11010111001010;     //141pi/512
  assign cos2[141]  =  14'b00110001010001;     //141pi/512
  assign sin2[142]  =  14'b11010110111011;     //142pi/512
  assign cos2[142]  =  14'b00110001000100;     //142pi/512
  assign sin2[143]  =  14'b11010110101011;     //143pi/512
  assign cos2[143]  =  14'b00110000110111;     //143pi/512
  assign sin2[144]  =  14'b11010110011100;     //144pi/512
  assign cos2[144]  =  14'b00110000101010;     //144pi/512
  assign sin2[145]  =  14'b11010110001101;     //145pi/512
  assign cos2[145]  =  14'b00110000011101;     //145pi/512
  assign sin2[146]  =  14'b11010101111101;     //146pi/512
  assign cos2[146]  =  14'b00110000010000;     //146pi/512
  assign sin2[147]  =  14'b11010101101110;     //147pi/512
  assign cos2[147]  =  14'b00110000000011;     //147pi/512
  assign sin2[148]  =  14'b11010101011111;     //148pi/512
  assign cos2[148]  =  14'b00101111110101;     //148pi/512
  assign sin2[149]  =  14'b11010101010000;     //149pi/512
  assign cos2[149]  =  14'b00101111101000;     //149pi/512
  assign sin2[150]  =  14'b11010101000001;     //150pi/512
  assign cos2[150]  =  14'b00101111011010;     //150pi/512
  assign sin2[151]  =  14'b11010100110010;     //151pi/512
  assign cos2[151]  =  14'b00101111001101;     //151pi/512
  assign sin2[152]  =  14'b11010100100100;     //152pi/512
  assign cos2[152]  =  14'b00101110111111;     //152pi/512
  assign sin2[153]  =  14'b11010100010101;     //153pi/512
  assign cos2[153]  =  14'b00101110110010;     //153pi/512
  assign sin2[154]  =  14'b11010100000110;     //154pi/512
  assign cos2[154]  =  14'b00101110100100;     //154pi/512
  assign sin2[155]  =  14'b11010011111000;     //155pi/512
  assign cos2[155]  =  14'b00101110010110;     //155pi/512
  assign sin2[156]  =  14'b11010011101001;     //156pi/512
  assign cos2[156]  =  14'b00101110001000;     //156pi/512
  assign sin2[157]  =  14'b11010011011011;     //157pi/512
  assign cos2[157]  =  14'b00101101111010;     //157pi/512
  assign sin2[158]  =  14'b11010011001100;     //158pi/512
  assign cos2[158]  =  14'b00101101101100;     //158pi/512
  assign sin2[159]  =  14'b11010010111110;     //159pi/512
  assign cos2[159]  =  14'b00101101011110;     //159pi/512
  assign sin2[160]  =  14'b11010010110000;     //160pi/512
  assign cos2[160]  =  14'b00101101010000;     //160pi/512
  assign sin2[161]  =  14'b11010010100010;     //161pi/512
  assign cos2[161]  =  14'b00101101000010;     //161pi/512
  assign sin2[162]  =  14'b11010010010011;     //162pi/512
  assign cos2[162]  =  14'b00101100110011;     //162pi/512
  assign sin2[163]  =  14'b11010010000101;     //163pi/512
  assign cos2[163]  =  14'b00101100100101;     //163pi/512
  assign sin2[164]  =  14'b11010001110111;     //164pi/512
  assign cos2[164]  =  14'b00101100010110;     //164pi/512
  assign sin2[165]  =  14'b11010001101001;     //165pi/512
  assign cos2[165]  =  14'b00101100001000;     //165pi/512
  assign sin2[166]  =  14'b11010001011100;     //166pi/512
  assign cos2[166]  =  14'b00101011111001;     //166pi/512
  assign sin2[167]  =  14'b11010001001110;     //167pi/512
  assign cos2[167]  =  14'b00101011101011;     //167pi/512
  assign sin2[168]  =  14'b11010001000000;     //168pi/512
  assign cos2[168]  =  14'b00101011011100;     //168pi/512
  assign sin2[169]  =  14'b11010000110011;     //169pi/512
  assign cos2[169]  =  14'b00101011001101;     //169pi/512
  assign sin2[170]  =  14'b11010000100101;     //170pi/512
  assign cos2[170]  =  14'b00101010111110;     //170pi/512
  assign sin2[171]  =  14'b11010000011000;     //171pi/512
  assign cos2[171]  =  14'b00101010101111;     //171pi/512
  assign sin2[172]  =  14'b11010000001010;     //172pi/512
  assign cos2[172]  =  14'b00101010100000;     //172pi/512
  assign sin2[173]  =  14'b11001111111101;     //173pi/512
  assign cos2[173]  =  14'b00101010010001;     //173pi/512
  assign sin2[174]  =  14'b11001111110000;     //174pi/512
  assign cos2[174]  =  14'b00101010000010;     //174pi/512
  assign sin2[175]  =  14'b11001111100010;     //175pi/512
  assign cos2[175]  =  14'b00101001110011;     //175pi/512
  assign sin2[176]  =  14'b11001111010101;     //176pi/512
  assign cos2[176]  =  14'b00101001100100;     //176pi/512
  assign sin2[177]  =  14'b11001111001000;     //177pi/512
  assign cos2[177]  =  14'b00101001010100;     //177pi/512
  assign sin2[178]  =  14'b11001110111011;     //178pi/512
  assign cos2[178]  =  14'b00101001000101;     //178pi/512
  assign sin2[179]  =  14'b11001110101111;     //179pi/512
  assign cos2[179]  =  14'b00101000110101;     //179pi/512
  assign sin2[180]  =  14'b11001110100010;     //180pi/512
  assign cos2[180]  =  14'b00101000100110;     //180pi/512
  assign sin2[181]  =  14'b11001110010101;     //181pi/512
  assign cos2[181]  =  14'b00101000010110;     //181pi/512
  assign sin2[182]  =  14'b11001110001000;     //182pi/512
  assign cos2[182]  =  14'b00101000000111;     //182pi/512
  assign sin2[183]  =  14'b11001101111100;     //183pi/512
  assign cos2[183]  =  14'b00100111110111;     //183pi/512
  assign sin2[184]  =  14'b11001101101111;     //184pi/512
  assign cos2[184]  =  14'b00100111100111;     //184pi/512
  assign sin2[185]  =  14'b11001101100011;     //185pi/512
  assign cos2[185]  =  14'b00100111010111;     //185pi/512
  assign sin2[186]  =  14'b11001101010111;     //186pi/512
  assign cos2[186]  =  14'b00100111001000;     //186pi/512
  assign sin2[187]  =  14'b11001101001010;     //187pi/512
  assign cos2[187]  =  14'b00100110111000;     //187pi/512
  assign sin2[188]  =  14'b11001100111110;     //188pi/512
  assign cos2[188]  =  14'b00100110101000;     //188pi/512
  assign sin2[189]  =  14'b11001100110010;     //189pi/512
  assign cos2[189]  =  14'b00100110011000;     //189pi/512
  assign sin2[190]  =  14'b11001100100110;     //190pi/512
  assign cos2[190]  =  14'b00100110000111;     //190pi/512
  assign sin2[191]  =  14'b11001100011010;     //191pi/512
  assign cos2[191]  =  14'b00100101110111;     //191pi/512
  assign sin2[192]  =  14'b11001100001110;     //192pi/512
  assign cos2[192]  =  14'b00100101100111;     //192pi/512
  assign sin2[193]  =  14'b11001100000010;     //193pi/512
  assign cos2[193]  =  14'b00100101010111;     //193pi/512
  assign sin2[194]  =  14'b11001011110111;     //194pi/512
  assign cos2[194]  =  14'b00100101000110;     //194pi/512
  assign sin2[195]  =  14'b11001011101011;     //195pi/512
  assign cos2[195]  =  14'b00100100110110;     //195pi/512
  assign sin2[196]  =  14'b11001011100000;     //196pi/512
  assign cos2[196]  =  14'b00100100100110;     //196pi/512
  assign sin2[197]  =  14'b11001011010100;     //197pi/512
  assign cos2[197]  =  14'b00100100010101;     //197pi/512
  assign sin2[198]  =  14'b11001011001001;     //198pi/512
  assign cos2[198]  =  14'b00100100000100;     //198pi/512
  assign sin2[199]  =  14'b11001010111110;     //199pi/512
  assign cos2[199]  =  14'b00100011110100;     //199pi/512
  assign sin2[200]  =  14'b11001010110010;     //200pi/512
  assign cos2[200]  =  14'b00100011100011;     //200pi/512
  assign sin2[201]  =  14'b11001010100111;     //201pi/512
  assign cos2[201]  =  14'b00100011010010;     //201pi/512
  assign sin2[202]  =  14'b11001010011100;     //202pi/512
  assign cos2[202]  =  14'b00100011000010;     //202pi/512
  assign sin2[203]  =  14'b11001010010001;     //203pi/512
  assign cos2[203]  =  14'b00100010110001;     //203pi/512
  assign sin2[204]  =  14'b11001010000110;     //204pi/512
  assign cos2[204]  =  14'b00100010100000;     //204pi/512
  assign sin2[205]  =  14'b11001001111011;     //205pi/512
  assign cos2[205]  =  14'b00100010001111;     //205pi/512
  assign sin2[206]  =  14'b11001001110001;     //206pi/512
  assign cos2[206]  =  14'b00100001111110;     //206pi/512
  assign sin2[207]  =  14'b11001001100110;     //207pi/512
  assign cos2[207]  =  14'b00100001101101;     //207pi/512
  assign sin2[208]  =  14'b11001001011100;     //208pi/512
  assign cos2[208]  =  14'b00100001011100;     //208pi/512
  assign sin2[209]  =  14'b11001001010001;     //209pi/512
  assign cos2[209]  =  14'b00100001001010;     //209pi/512
  assign sin2[210]  =  14'b11001001000111;     //210pi/512
  assign cos2[210]  =  14'b00100000111001;     //210pi/512
  assign sin2[211]  =  14'b11001000111100;     //211pi/512
  assign cos2[211]  =  14'b00100000101000;     //211pi/512
  assign sin2[212]  =  14'b11001000110010;     //212pi/512
  assign cos2[212]  =  14'b00100000010111;     //212pi/512
  assign sin2[213]  =  14'b11001000101000;     //213pi/512
  assign cos2[213]  =  14'b00100000000101;     //213pi/512
  assign sin2[214]  =  14'b11001000011110;     //214pi/512
  assign cos2[214]  =  14'b00011111110100;     //214pi/512
  assign sin2[215]  =  14'b11001000010100;     //215pi/512
  assign cos2[215]  =  14'b00011111100010;     //215pi/512
  assign sin2[216]  =  14'b11001000001010;     //216pi/512
  assign cos2[216]  =  14'b00011111010001;     //216pi/512
  assign sin2[217]  =  14'b11001000000000;     //217pi/512
  assign cos2[217]  =  14'b00011110111111;     //217pi/512
  assign sin2[218]  =  14'b11000111110111;     //218pi/512
  assign cos2[218]  =  14'b00011110101110;     //218pi/512
  assign sin2[219]  =  14'b11000111101101;     //219pi/512
  assign cos2[219]  =  14'b00011110011100;     //219pi/512
  assign sin2[220]  =  14'b11000111100100;     //220pi/512
  assign cos2[220]  =  14'b00011110001010;     //220pi/512
  assign sin2[221]  =  14'b11000111011010;     //221pi/512
  assign cos2[221]  =  14'b00011101111001;     //221pi/512
  assign sin2[222]  =  14'b11000111010001;     //222pi/512
  assign cos2[222]  =  14'b00011101100111;     //222pi/512
  assign sin2[223]  =  14'b11000111001000;     //223pi/512
  assign cos2[223]  =  14'b00011101010101;     //223pi/512
  assign sin2[224]  =  14'b11000110111110;     //224pi/512
  assign cos2[224]  =  14'b00011101000011;     //224pi/512
  assign sin2[225]  =  14'b11000110110101;     //225pi/512
  assign cos2[225]  =  14'b00011100110001;     //225pi/512
  assign sin2[226]  =  14'b11000110101100;     //226pi/512
  assign cos2[226]  =  14'b00011100011111;     //226pi/512
  assign sin2[227]  =  14'b11000110100011;     //227pi/512
  assign cos2[227]  =  14'b00011100001101;     //227pi/512
  assign sin2[228]  =  14'b11000110011011;     //228pi/512
  assign cos2[228]  =  14'b00011011111011;     //228pi/512
  assign sin2[229]  =  14'b11000110010010;     //229pi/512
  assign cos2[229]  =  14'b00011011101001;     //229pi/512
  assign sin2[230]  =  14'b11000110001001;     //230pi/512
  assign cos2[230]  =  14'b00011011010111;     //230pi/512
  assign sin2[231]  =  14'b11000110000001;     //231pi/512
  assign cos2[231]  =  14'b00011011000101;     //231pi/512
  assign sin2[232]  =  14'b11000101111000;     //232pi/512
  assign cos2[232]  =  14'b00011010110010;     //232pi/512
  assign sin2[233]  =  14'b11000101110000;     //233pi/512
  assign cos2[233]  =  14'b00011010100000;     //233pi/512
  assign sin2[234]  =  14'b11000101101000;     //234pi/512
  assign cos2[234]  =  14'b00011010001110;     //234pi/512
  assign sin2[235]  =  14'b11000101011111;     //235pi/512
  assign cos2[235]  =  14'b00011001111011;     //235pi/512
  assign sin2[236]  =  14'b11000101010111;     //236pi/512
  assign cos2[236]  =  14'b00011001101001;     //236pi/512
  assign sin2[237]  =  14'b11000101001111;     //237pi/512
  assign cos2[237]  =  14'b00011001010111;     //237pi/512
  assign sin2[238]  =  14'b11000101000111;     //238pi/512
  assign cos2[238]  =  14'b00011001000100;     //238pi/512
  assign sin2[239]  =  14'b11000101000000;     //239pi/512
  assign cos2[239]  =  14'b00011000110010;     //239pi/512
  assign sin2[240]  =  14'b11000100111000;     //240pi/512
  assign cos2[240]  =  14'b00011000011111;     //240pi/512
  assign sin2[241]  =  14'b11000100110000;     //241pi/512
  assign cos2[241]  =  14'b00011000001100;     //241pi/512
  assign sin2[242]  =  14'b11000100101001;     //242pi/512
  assign cos2[242]  =  14'b00010111111010;     //242pi/512
  assign sin2[243]  =  14'b11000100100001;     //243pi/512
  assign cos2[243]  =  14'b00010111100111;     //243pi/512
  assign sin2[244]  =  14'b11000100011010;     //244pi/512
  assign cos2[244]  =  14'b00010111010100;     //244pi/512
  assign sin2[245]  =  14'b11000100010010;     //245pi/512
  assign cos2[245]  =  14'b00010111000010;     //245pi/512
  assign sin2[246]  =  14'b11000100001011;     //246pi/512
  assign cos2[246]  =  14'b00010110101111;     //246pi/512
  assign sin2[247]  =  14'b11000100000100;     //247pi/512
  assign cos2[247]  =  14'b00010110011100;     //247pi/512
  assign sin2[248]  =  14'b11000011111101;     //248pi/512
  assign cos2[248]  =  14'b00010110001001;     //248pi/512
  assign sin2[249]  =  14'b11000011110110;     //249pi/512
  assign cos2[249]  =  14'b00010101110110;     //249pi/512
  assign sin2[250]  =  14'b11000011101111;     //250pi/512
  assign cos2[250]  =  14'b00010101100011;     //250pi/512
  assign sin2[251]  =  14'b11000011101001;     //251pi/512
  assign cos2[251]  =  14'b00010101010000;     //251pi/512
  assign sin2[252]  =  14'b11000011100010;     //252pi/512
  assign cos2[252]  =  14'b00010100111101;     //252pi/512
  assign sin2[253]  =  14'b11000011011100;     //253pi/512
  assign cos2[253]  =  14'b00010100101010;     //253pi/512
  assign sin2[254]  =  14'b11000011010101;     //254pi/512
  assign cos2[254]  =  14'b00010100010111;     //254pi/512
  assign sin2[255]  =  14'b11000011001111;     //255pi/512
  assign cos2[255]  =  14'b00010100000100;     //255pi/512
  assign sin2[256]  =  14'b11000011001000;     //256pi/512
  assign cos2[256]  =  14'b00010011110001;     //256pi/512
  assign sin2[257]  =  14'b11000011000010;     //257pi/512
  assign cos2[257]  =  14'b00010011011110;     //257pi/512
  assign sin2[258]  =  14'b11000010111100;     //258pi/512
  assign cos2[258]  =  14'b00010011001011;     //258pi/512
  assign sin2[259]  =  14'b11000010110110;     //259pi/512
  assign cos2[259]  =  14'b00010010111000;     //259pi/512
  assign sin2[260]  =  14'b11000010110000;     //260pi/512
  assign cos2[260]  =  14'b00010010100101;     //260pi/512
  assign sin2[261]  =  14'b11000010101011;     //261pi/512
  assign cos2[261]  =  14'b00010010010001;     //261pi/512
  assign sin2[262]  =  14'b11000010100101;     //262pi/512
  assign cos2[262]  =  14'b00010001111110;     //262pi/512
  assign sin2[263]  =  14'b11000010011111;     //263pi/512
  assign cos2[263]  =  14'b00010001101011;     //263pi/512
  assign sin2[264]  =  14'b11000010011010;     //264pi/512
  assign cos2[264]  =  14'b00010001010111;     //264pi/512
  assign sin2[265]  =  14'b11000010010100;     //265pi/512
  assign cos2[265]  =  14'b00010001000100;     //265pi/512
  assign sin2[266]  =  14'b11000010001111;     //266pi/512
  assign cos2[266]  =  14'b00010000110001;     //266pi/512
  assign sin2[267]  =  14'b11000010001010;     //267pi/512
  assign cos2[267]  =  14'b00010000011101;     //267pi/512
  assign sin2[268]  =  14'b11000010000101;     //268pi/512
  assign cos2[268]  =  14'b00010000001010;     //268pi/512
  assign sin2[269]  =  14'b11000010000000;     //269pi/512
  assign cos2[269]  =  14'b00001111110110;     //269pi/512
  assign sin2[270]  =  14'b11000001111011;     //270pi/512
  assign cos2[270]  =  14'b00001111100011;     //270pi/512
  assign sin2[271]  =  14'b11000001110110;     //271pi/512
  assign cos2[271]  =  14'b00001111001111;     //271pi/512
  assign sin2[272]  =  14'b11000001110001;     //272pi/512
  assign cos2[272]  =  14'b00001110111100;     //272pi/512
  assign sin2[273]  =  14'b11000001101101;     //273pi/512
  assign cos2[273]  =  14'b00001110101000;     //273pi/512
  assign sin2[274]  =  14'b11000001101000;     //274pi/512
  assign cos2[274]  =  14'b00001110010101;     //274pi/512
  assign sin2[275]  =  14'b11000001100100;     //275pi/512
  assign cos2[275]  =  14'b00001110000001;     //275pi/512
  assign sin2[276]  =  14'b11000001011111;     //276pi/512
  assign cos2[276]  =  14'b00001101101101;     //276pi/512
  assign sin2[277]  =  14'b11000001011011;     //277pi/512
  assign cos2[277]  =  14'b00001101011010;     //277pi/512
  assign sin2[278]  =  14'b11000001010111;     //278pi/512
  assign cos2[278]  =  14'b00001101000110;     //278pi/512
  assign sin2[279]  =  14'b11000001010011;     //279pi/512
  assign cos2[279]  =  14'b00001100110010;     //279pi/512
  assign sin2[280]  =  14'b11000001001111;     //280pi/512
  assign cos2[280]  =  14'b00001100011111;     //280pi/512
  assign sin2[281]  =  14'b11000001001011;     //281pi/512
  assign cos2[281]  =  14'b00001100001011;     //281pi/512
  assign sin2[282]  =  14'b11000001000111;     //282pi/512
  assign cos2[282]  =  14'b00001011110111;     //282pi/512
  assign sin2[283]  =  14'b11000001000011;     //283pi/512
  assign cos2[283]  =  14'b00001011100011;     //283pi/512
  assign sin2[284]  =  14'b11000001000000;     //284pi/512
  assign cos2[284]  =  14'b00001011010000;     //284pi/512
  assign sin2[285]  =  14'b11000000111100;     //285pi/512
  assign cos2[285]  =  14'b00001010111100;     //285pi/512
  assign sin2[286]  =  14'b11000000111001;     //286pi/512
  assign cos2[286]  =  14'b00001010101000;     //286pi/512
  assign sin2[287]  =  14'b11000000110110;     //287pi/512
  assign cos2[287]  =  14'b00001010010100;     //287pi/512
  assign sin2[288]  =  14'b11000000110010;     //288pi/512
  assign cos2[288]  =  14'b00001010000000;     //288pi/512
  assign sin2[289]  =  14'b11000000101111;     //289pi/512
  assign cos2[289]  =  14'b00001001101100;     //289pi/512
  assign sin2[290]  =  14'b11000000101100;     //290pi/512
  assign cos2[290]  =  14'b00001001011001;     //290pi/512
  assign sin2[291]  =  14'b11000000101001;     //291pi/512
  assign cos2[291]  =  14'b00001001000101;     //291pi/512
  assign sin2[292]  =  14'b11000000100111;     //292pi/512
  assign cos2[292]  =  14'b00001000110001;     //292pi/512
  assign sin2[293]  =  14'b11000000100100;     //293pi/512
  assign cos2[293]  =  14'b00001000011101;     //293pi/512
  assign sin2[294]  =  14'b11000000100001;     //294pi/512
  assign cos2[294]  =  14'b00001000001001;     //294pi/512
  assign sin2[295]  =  14'b11000000011111;     //295pi/512
  assign cos2[295]  =  14'b00000111110101;     //295pi/512
  assign sin2[296]  =  14'b11000000011100;     //296pi/512
  assign cos2[296]  =  14'b00000111100001;     //296pi/512
  assign sin2[297]  =  14'b11000000011010;     //297pi/512
  assign cos2[297]  =  14'b00000111001101;     //297pi/512
  assign sin2[298]  =  14'b11000000011000;     //298pi/512
  assign cos2[298]  =  14'b00000110111001;     //298pi/512
  assign sin2[299]  =  14'b11000000010110;     //299pi/512
  assign cos2[299]  =  14'b00000110100101;     //299pi/512
  assign sin2[300]  =  14'b11000000010100;     //300pi/512
  assign cos2[300]  =  14'b00000110010001;     //300pi/512
  assign sin2[301]  =  14'b11000000010010;     //301pi/512
  assign cos2[301]  =  14'b00000101111101;     //301pi/512
  assign sin2[302]  =  14'b11000000010000;     //302pi/512
  assign cos2[302]  =  14'b00000101101001;     //302pi/512
  assign sin2[303]  =  14'b11000000001110;     //303pi/512
  assign cos2[303]  =  14'b00000101010101;     //303pi/512
  assign sin2[304]  =  14'b11000000001101;     //304pi/512
  assign cos2[304]  =  14'b00000101000001;     //304pi/512
  assign sin2[305]  =  14'b11000000001011;     //305pi/512
  assign cos2[305]  =  14'b00000100101101;     //305pi/512
  assign sin2[306]  =  14'b11000000001010;     //306pi/512
  assign cos2[306]  =  14'b00000100011001;     //306pi/512
  assign sin2[307]  =  14'b11000000001000;     //307pi/512
  assign cos2[307]  =  14'b00000100000101;     //307pi/512
  assign sin2[308]  =  14'b11000000000111;     //308pi/512
  assign cos2[308]  =  14'b00000011110001;     //308pi/512
  assign sin2[309]  =  14'b11000000000110;     //309pi/512
  assign cos2[309]  =  14'b00000011011101;     //309pi/512
  assign sin2[310]  =  14'b11000000000101;     //310pi/512
  assign cos2[310]  =  14'b00000011001000;     //310pi/512
  assign sin2[311]  =  14'b11000000000100;     //311pi/512
  assign cos2[311]  =  14'b00000010110100;     //311pi/512
  assign sin2[312]  =  14'b11000000000011;     //312pi/512
  assign cos2[312]  =  14'b00000010100000;     //312pi/512
  assign sin2[313]  =  14'b11000000000010;     //313pi/512
  assign cos2[313]  =  14'b00000010001100;     //313pi/512
  assign sin2[314]  =  14'b11000000000010;     //314pi/512
  assign cos2[314]  =  14'b00000001111000;     //314pi/512
  assign sin2[315]  =  14'b11000000000001;     //315pi/512
  assign cos2[315]  =  14'b00000001100100;     //315pi/512
  assign sin2[316]  =  14'b11000000000001;     //316pi/512
  assign cos2[316]  =  14'b00000001010000;     //316pi/512
  assign sin2[317]  =  14'b11000000000000;     //317pi/512
  assign cos2[317]  =  14'b00000000111100;     //317pi/512
  assign sin2[318]  =  14'b11000000000000;     //318pi/512
  assign cos2[318]  =  14'b00000000101000;     //318pi/512
  assign sin2[319]  =  14'b11000000000000;     //319pi/512
  assign cos2[319]  =  14'b00000000010100;     //319pi/512
  assign sin2[320]  =  14'b11000000000000;     //320pi/512
  assign cos2[320]  =  14'b00000000000000;     //320pi/512
  assign sin2[321]  =  14'b11000000000000;     //321pi/512
  assign cos2[321]  =  14'b11111111101100;     //321pi/512
  assign sin2[322]  =  14'b11000000000000;     //322pi/512
  assign cos2[322]  =  14'b11111111011000;     //322pi/512
  assign sin2[323]  =  14'b11000000000000;     //323pi/512
  assign cos2[323]  =  14'b11111111000100;     //323pi/512
  assign sin2[324]  =  14'b11000000000001;     //324pi/512
  assign cos2[324]  =  14'b11111110110000;     //324pi/512
  assign sin2[325]  =  14'b11000000000001;     //325pi/512
  assign cos2[325]  =  14'b11111110011011;     //325pi/512
  assign sin2[326]  =  14'b11000000000010;     //326pi/512
  assign cos2[326]  =  14'b11111110000111;     //326pi/512
  assign sin2[327]  =  14'b11000000000010;     //327pi/512
  assign cos2[327]  =  14'b11111101110011;     //327pi/512
  assign sin2[328]  =  14'b11000000000011;     //328pi/512
  assign cos2[328]  =  14'b11111101011111;     //328pi/512
  assign sin2[329]  =  14'b11000000000100;     //329pi/512
  assign cos2[329]  =  14'b11111101001011;     //329pi/512
  assign sin2[330]  =  14'b11000000000101;     //330pi/512
  assign cos2[330]  =  14'b11111100110111;     //330pi/512
  assign sin2[331]  =  14'b11000000000110;     //331pi/512
  assign cos2[331]  =  14'b11111100100011;     //331pi/512
  assign sin2[332]  =  14'b11000000000111;     //332pi/512
  assign cos2[332]  =  14'b11111100001111;     //332pi/512
  assign sin2[333]  =  14'b11000000001000;     //333pi/512
  assign cos2[333]  =  14'b11111011111011;     //333pi/512
  assign sin2[334]  =  14'b11000000001010;     //334pi/512
  assign cos2[334]  =  14'b11111011100111;     //334pi/512
  assign sin2[335]  =  14'b11000000001011;     //335pi/512
  assign cos2[335]  =  14'b11111011010011;     //335pi/512
  assign sin2[336]  =  14'b11000000001101;     //336pi/512
  assign cos2[336]  =  14'b11111010111111;     //336pi/512
  assign sin2[337]  =  14'b11000000001110;     //337pi/512
  assign cos2[337]  =  14'b11111010101011;     //337pi/512
  assign sin2[338]  =  14'b11000000010000;     //338pi/512
  assign cos2[338]  =  14'b11111010010111;     //338pi/512
  assign sin2[339]  =  14'b11000000010010;     //339pi/512
  assign cos2[339]  =  14'b11111010000011;     //339pi/512
  assign sin2[340]  =  14'b11000000010100;     //340pi/512
  assign cos2[340]  =  14'b11111001101111;     //340pi/512
  assign sin2[341]  =  14'b11000000010110;     //341pi/512
  assign cos2[341]  =  14'b11111001011011;     //341pi/512
  assign sin2[342]  =  14'b11000000011000;     //342pi/512
  assign cos2[342]  =  14'b11111001000111;     //342pi/512
  assign sin2[343]  =  14'b11000000011010;     //343pi/512
  assign cos2[343]  =  14'b11111000110011;     //343pi/512
  assign sin2[344]  =  14'b11000000011100;     //344pi/512
  assign cos2[344]  =  14'b11111000011111;     //344pi/512
  assign sin2[345]  =  14'b11000000011111;     //345pi/512
  assign cos2[345]  =  14'b11111000001011;     //345pi/512
  assign sin2[346]  =  14'b11000000100001;     //346pi/512
  assign cos2[346]  =  14'b11110111110111;     //346pi/512
  assign sin2[347]  =  14'b11000000100100;     //347pi/512
  assign cos2[347]  =  14'b11110111100011;     //347pi/512
  assign sin2[348]  =  14'b11000000100111;     //348pi/512
  assign cos2[348]  =  14'b11110111001111;     //348pi/512
  assign sin2[349]  =  14'b11000000101001;     //349pi/512
  assign cos2[349]  =  14'b11110110111011;     //349pi/512
  assign sin2[350]  =  14'b11000000101100;     //350pi/512
  assign cos2[350]  =  14'b11110110100111;     //350pi/512
  assign sin2[351]  =  14'b11000000101111;     //351pi/512
  assign cos2[351]  =  14'b11110110010011;     //351pi/512
  assign sin2[352]  =  14'b11000000110010;     //352pi/512
  assign cos2[352]  =  14'b11110101111111;     //352pi/512
  assign sin2[353]  =  14'b11000000110110;     //353pi/512
  assign cos2[353]  =  14'b11110101101011;     //353pi/512
  assign sin2[354]  =  14'b11000000111001;     //354pi/512
  assign cos2[354]  =  14'b11110101011000;     //354pi/512
  assign sin2[355]  =  14'b11000000111100;     //355pi/512
  assign cos2[355]  =  14'b11110101000100;     //355pi/512
  assign sin2[356]  =  14'b11000001000000;     //356pi/512
  assign cos2[356]  =  14'b11110100110000;     //356pi/512
  assign sin2[357]  =  14'b11000001000011;     //357pi/512
  assign cos2[357]  =  14'b11110100011100;     //357pi/512
  assign sin2[358]  =  14'b11000001000111;     //358pi/512
  assign cos2[358]  =  14'b11110100001000;     //358pi/512
  assign sin2[359]  =  14'b11000001001011;     //359pi/512
  assign cos2[359]  =  14'b11110011110101;     //359pi/512
  assign sin2[360]  =  14'b11000001001111;     //360pi/512
  assign cos2[360]  =  14'b11110011100001;     //360pi/512
  assign sin2[361]  =  14'b11000001010011;     //361pi/512
  assign cos2[361]  =  14'b11110011001101;     //361pi/512
  assign sin2[362]  =  14'b11000001010111;     //362pi/512
  assign cos2[362]  =  14'b11110010111010;     //362pi/512
  assign sin2[363]  =  14'b11000001011011;     //363pi/512
  assign cos2[363]  =  14'b11110010100110;     //363pi/512
  assign sin2[364]  =  14'b11000001011111;     //364pi/512
  assign cos2[364]  =  14'b11110010010010;     //364pi/512
  assign sin2[365]  =  14'b11000001100100;     //365pi/512
  assign cos2[365]  =  14'b11110001111111;     //365pi/512
  assign sin2[366]  =  14'b11000001101000;     //366pi/512
  assign cos2[366]  =  14'b11110001101011;     //366pi/512
  assign sin2[367]  =  14'b11000001101101;     //367pi/512
  assign cos2[367]  =  14'b11110001010111;     //367pi/512
  assign sin2[368]  =  14'b11000001110001;     //368pi/512
  assign cos2[368]  =  14'b11110001000100;     //368pi/512
  assign sin2[369]  =  14'b11000001110110;     //369pi/512
  assign cos2[369]  =  14'b11110000110000;     //369pi/512
  assign sin2[370]  =  14'b11000001111011;     //370pi/512
  assign cos2[370]  =  14'b11110000011101;     //370pi/512
  assign sin2[371]  =  14'b11000010000000;     //371pi/512
  assign cos2[371]  =  14'b11110000001001;     //371pi/512
  assign sin2[372]  =  14'b11000010000101;     //372pi/512
  assign cos2[372]  =  14'b11101111110110;     //372pi/512
  assign sin2[373]  =  14'b11000010001010;     //373pi/512
  assign cos2[373]  =  14'b11101111100010;     //373pi/512
  assign sin2[374]  =  14'b11000010001111;     //374pi/512
  assign cos2[374]  =  14'b11101111001111;     //374pi/512
  assign sin2[375]  =  14'b11000010010100;     //375pi/512
  assign cos2[375]  =  14'b11101110111100;     //375pi/512
  assign sin2[376]  =  14'b11000010011010;     //376pi/512
  assign cos2[376]  =  14'b11101110101000;     //376pi/512
  assign sin2[377]  =  14'b11000010011111;     //377pi/512
  assign cos2[377]  =  14'b11101110010101;     //377pi/512
  assign sin2[378]  =  14'b11000010100101;     //378pi/512
  assign cos2[378]  =  14'b11101110000010;     //378pi/512
  assign sin2[379]  =  14'b11000010101011;     //379pi/512
  assign cos2[379]  =  14'b11101101101110;     //379pi/512
  assign sin2[380]  =  14'b11000010110000;     //380pi/512
  assign cos2[380]  =  14'b11101101011011;     //380pi/512
  assign sin2[381]  =  14'b11000010110110;     //381pi/512
  assign cos2[381]  =  14'b11101101001000;     //381pi/512
  assign sin2[382]  =  14'b11000010111100;     //382pi/512
  assign cos2[382]  =  14'b11101100110101;     //382pi/512
  assign sin2[383]  =  14'b11000011000010;     //383pi/512
  assign cos2[383]  =  14'b11101100100001;     //383pi/512
  assign sin2[384]  =  14'b11000011001000;     //384pi/512
  assign cos2[384]  =  14'b11101100001110;     //384pi/512
  assign sin2[385]  =  14'b11000011001111;     //385pi/512
  assign cos2[385]  =  14'b11101011111011;     //385pi/512
  assign sin2[386]  =  14'b11000011010101;     //386pi/512
  assign cos2[386]  =  14'b11101011101000;     //386pi/512
  assign sin2[387]  =  14'b11000011011100;     //387pi/512
  assign cos2[387]  =  14'b11101011010101;     //387pi/512
  assign sin2[388]  =  14'b11000011100010;     //388pi/512
  assign cos2[388]  =  14'b11101011000010;     //388pi/512
  assign sin2[389]  =  14'b11000011101001;     //389pi/512
  assign cos2[389]  =  14'b11101010101111;     //389pi/512
  assign sin2[390]  =  14'b11000011101111;     //390pi/512
  assign cos2[390]  =  14'b11101010011100;     //390pi/512
  assign sin2[391]  =  14'b11000011110110;     //391pi/512
  assign cos2[391]  =  14'b11101010001001;     //391pi/512
  assign sin2[392]  =  14'b11000011111101;     //392pi/512
  assign cos2[392]  =  14'b11101001110110;     //392pi/512
  assign sin2[393]  =  14'b11000100000100;     //393pi/512
  assign cos2[393]  =  14'b11101001100011;     //393pi/512
  assign sin2[394]  =  14'b11000100001011;     //394pi/512
  assign cos2[394]  =  14'b11101001010001;     //394pi/512
  assign sin2[395]  =  14'b11000100010010;     //395pi/512
  assign cos2[395]  =  14'b11101000111110;     //395pi/512
  assign sin2[396]  =  14'b11000100011010;     //396pi/512
  assign cos2[396]  =  14'b11101000101011;     //396pi/512
  assign sin2[397]  =  14'b11000100100001;     //397pi/512
  assign cos2[397]  =  14'b11101000011000;     //397pi/512
  assign sin2[398]  =  14'b11000100101001;     //398pi/512
  assign cos2[398]  =  14'b11101000000110;     //398pi/512
  assign sin2[399]  =  14'b11000100110000;     //399pi/512
  assign cos2[399]  =  14'b11100111110011;     //399pi/512
  assign sin2[400]  =  14'b11000100111000;     //400pi/512
  assign cos2[400]  =  14'b11100111100001;     //400pi/512
  assign sin2[401]  =  14'b11000101000000;     //401pi/512
  assign cos2[401]  =  14'b11100111001110;     //401pi/512
  assign sin2[402]  =  14'b11000101000111;     //402pi/512
  assign cos2[402]  =  14'b11100110111011;     //402pi/512
  assign sin2[403]  =  14'b11000101001111;     //403pi/512
  assign cos2[403]  =  14'b11100110101001;     //403pi/512
  assign sin2[404]  =  14'b11000101010111;     //404pi/512
  assign cos2[404]  =  14'b11100110010111;     //404pi/512
  assign sin2[405]  =  14'b11000101011111;     //405pi/512
  assign cos2[405]  =  14'b11100110000100;     //405pi/512
  assign sin2[406]  =  14'b11000101101000;     //406pi/512
  assign cos2[406]  =  14'b11100101110010;     //406pi/512
  assign sin2[407]  =  14'b11000101110000;     //407pi/512
  assign cos2[407]  =  14'b11100101011111;     //407pi/512
  assign sin2[408]  =  14'b11000101111000;     //408pi/512
  assign cos2[408]  =  14'b11100101001101;     //408pi/512
  assign sin2[409]  =  14'b11000110000001;     //409pi/512
  assign cos2[409]  =  14'b11100100111011;     //409pi/512
  assign sin2[410]  =  14'b11000110001001;     //410pi/512
  assign cos2[410]  =  14'b11100100101001;     //410pi/512
  assign sin2[411]  =  14'b11000110010010;     //411pi/512
  assign cos2[411]  =  14'b11100100010111;     //411pi/512
  assign sin2[412]  =  14'b11000110011011;     //412pi/512
  assign cos2[412]  =  14'b11100100000100;     //412pi/512
  assign sin2[413]  =  14'b11000110100011;     //413pi/512
  assign cos2[413]  =  14'b11100011110010;     //413pi/512
  assign sin2[414]  =  14'b11000110101100;     //414pi/512
  assign cos2[414]  =  14'b11100011100000;     //414pi/512
  assign sin2[415]  =  14'b11000110110101;     //415pi/512
  assign cos2[415]  =  14'b11100011001110;     //415pi/512
  assign sin2[416]  =  14'b11000110111110;     //416pi/512
  assign cos2[416]  =  14'b11100010111100;     //416pi/512
  assign sin2[417]  =  14'b11000111001000;     //417pi/512
  assign cos2[417]  =  14'b11100010101011;     //417pi/512
  assign sin2[418]  =  14'b11000111010001;     //418pi/512
  assign cos2[418]  =  14'b11100010011001;     //418pi/512
  assign sin2[419]  =  14'b11000111011010;     //419pi/512
  assign cos2[419]  =  14'b11100010000111;     //419pi/512
  assign sin2[420]  =  14'b11000111100100;     //420pi/512
  assign cos2[420]  =  14'b11100001110101;     //420pi/512
  assign sin2[421]  =  14'b11000111101101;     //421pi/512
  assign cos2[421]  =  14'b11100001100011;     //421pi/512
  assign sin2[422]  =  14'b11000111110111;     //422pi/512
  assign cos2[422]  =  14'b11100001010010;     //422pi/512
  assign sin2[423]  =  14'b11001000000000;     //423pi/512
  assign cos2[423]  =  14'b11100001000000;     //423pi/512
  assign sin2[424]  =  14'b11001000001010;     //424pi/512
  assign cos2[424]  =  14'b11100000101111;     //424pi/512
  assign sin2[425]  =  14'b11001000010100;     //425pi/512
  assign cos2[425]  =  14'b11100000011101;     //425pi/512
  assign sin2[426]  =  14'b11001000011110;     //426pi/512
  assign cos2[426]  =  14'b11100000001100;     //426pi/512
  assign sin2[427]  =  14'b11001000101000;     //427pi/512
  assign cos2[427]  =  14'b11011111111010;     //427pi/512
  assign sin2[428]  =  14'b11001000110010;     //428pi/512
  assign cos2[428]  =  14'b11011111101001;     //428pi/512
  assign sin2[429]  =  14'b11001000111100;     //429pi/512
  assign cos2[429]  =  14'b11011111011000;     //429pi/512
  assign sin2[430]  =  14'b11001001000111;     //430pi/512
  assign cos2[430]  =  14'b11011111000110;     //430pi/512
  assign sin2[431]  =  14'b11001001010001;     //431pi/512
  assign cos2[431]  =  14'b11011110110101;     //431pi/512
  assign sin2[432]  =  14'b11001001011100;     //432pi/512
  assign cos2[432]  =  14'b11011110100100;     //432pi/512
  assign sin2[433]  =  14'b11001001100110;     //433pi/512
  assign cos2[433]  =  14'b11011110010011;     //433pi/512
  assign sin2[434]  =  14'b11001001110001;     //434pi/512
  assign cos2[434]  =  14'b11011110000010;     //434pi/512
  assign sin2[435]  =  14'b11001001111011;     //435pi/512
  assign cos2[435]  =  14'b11011101110001;     //435pi/512
  assign sin2[436]  =  14'b11001010000110;     //436pi/512
  assign cos2[436]  =  14'b11011101100000;     //436pi/512
  assign sin2[437]  =  14'b11001010010001;     //437pi/512
  assign cos2[437]  =  14'b11011101001111;     //437pi/512
  assign sin2[438]  =  14'b11001010011100;     //438pi/512
  assign cos2[438]  =  14'b11011100111110;     //438pi/512
  assign sin2[439]  =  14'b11001010100111;     //439pi/512
  assign cos2[439]  =  14'b11011100101101;     //439pi/512
  assign sin2[440]  =  14'b11001010110010;     //440pi/512
  assign cos2[440]  =  14'b11011100011100;     //440pi/512
  assign sin2[441]  =  14'b11001010111110;     //441pi/512
  assign cos2[441]  =  14'b11011100001100;     //441pi/512
  assign sin2[442]  =  14'b11001011001001;     //442pi/512
  assign cos2[442]  =  14'b11011011111011;     //442pi/512
  assign sin2[443]  =  14'b11001011010100;     //443pi/512
  assign cos2[443]  =  14'b11011011101010;     //443pi/512
  assign sin2[444]  =  14'b11001011100000;     //444pi/512
  assign cos2[444]  =  14'b11011011011010;     //444pi/512
  assign sin2[445]  =  14'b11001011101011;     //445pi/512
  assign cos2[445]  =  14'b11011011001001;     //445pi/512
  assign sin2[446]  =  14'b11001011110111;     //446pi/512
  assign cos2[446]  =  14'b11011010111001;     //446pi/512
  assign sin2[447]  =  14'b11001100000010;     //447pi/512
  assign cos2[447]  =  14'b11011010101001;     //447pi/512
  assign sin2[448]  =  14'b11001100001110;     //448pi/512
  assign cos2[448]  =  14'b11011010011000;     //448pi/512
  assign sin2[449]  =  14'b11001100011010;     //449pi/512
  assign cos2[449]  =  14'b11011010001000;     //449pi/512
  assign sin2[450]  =  14'b11001100100110;     //450pi/512
  assign cos2[450]  =  14'b11011001111000;     //450pi/512
  assign sin2[451]  =  14'b11001100110010;     //451pi/512
  assign cos2[451]  =  14'b11011001101000;     //451pi/512
  assign sin2[452]  =  14'b11001100111110;     //452pi/512
  assign cos2[452]  =  14'b11011001011000;     //452pi/512
  assign sin2[453]  =  14'b11001101001010;     //453pi/512
  assign cos2[453]  =  14'b11011001001000;     //453pi/512
  assign sin2[454]  =  14'b11001101010111;     //454pi/512
  assign cos2[454]  =  14'b11011000111000;     //454pi/512
  assign sin2[455]  =  14'b11001101100011;     //455pi/512
  assign cos2[455]  =  14'b11011000101000;     //455pi/512
  assign sin2[456]  =  14'b11001101101111;     //456pi/512
  assign cos2[456]  =  14'b11011000011000;     //456pi/512
  assign sin2[457]  =  14'b11001101111100;     //457pi/512
  assign cos2[457]  =  14'b11011000001000;     //457pi/512
  assign sin2[458]  =  14'b11001110001000;     //458pi/512
  assign cos2[458]  =  14'b11010111111001;     //458pi/512
  assign sin2[459]  =  14'b11001110010101;     //459pi/512
  assign cos2[459]  =  14'b11010111101001;     //459pi/512
  assign sin2[460]  =  14'b11001110100010;     //460pi/512
  assign cos2[460]  =  14'b11010111011010;     //460pi/512
  assign sin2[461]  =  14'b11001110101111;     //461pi/512
  assign cos2[461]  =  14'b11010111001010;     //461pi/512
  assign sin2[462]  =  14'b11001110111011;     //462pi/512
  assign cos2[462]  =  14'b11010110111011;     //462pi/512
  assign sin2[463]  =  14'b11001111001000;     //463pi/512
  assign cos2[463]  =  14'b11010110101011;     //463pi/512
  assign sin2[464]  =  14'b11001111010101;     //464pi/512
  assign cos2[464]  =  14'b11010110011100;     //464pi/512
  assign sin2[465]  =  14'b11001111100010;     //465pi/512
  assign cos2[465]  =  14'b11010110001101;     //465pi/512
  assign sin2[466]  =  14'b11001111110000;     //466pi/512
  assign cos2[466]  =  14'b11010101111101;     //466pi/512
  assign sin2[467]  =  14'b11001111111101;     //467pi/512
  assign cos2[467]  =  14'b11010101101110;     //467pi/512
  assign sin2[468]  =  14'b11010000001010;     //468pi/512
  assign cos2[468]  =  14'b11010101011111;     //468pi/512
  assign sin2[469]  =  14'b11010000011000;     //469pi/512
  assign cos2[469]  =  14'b11010101010000;     //469pi/512
  assign sin2[470]  =  14'b11010000100101;     //470pi/512
  assign cos2[470]  =  14'b11010101000001;     //470pi/512
  assign sin2[471]  =  14'b11010000110011;     //471pi/512
  assign cos2[471]  =  14'b11010100110010;     //471pi/512
  assign sin2[472]  =  14'b11010001000000;     //472pi/512
  assign cos2[472]  =  14'b11010100100100;     //472pi/512
  assign sin2[473]  =  14'b11010001001110;     //473pi/512
  assign cos2[473]  =  14'b11010100010101;     //473pi/512
  assign sin2[474]  =  14'b11010001011100;     //474pi/512
  assign cos2[474]  =  14'b11010100000110;     //474pi/512
  assign sin2[475]  =  14'b11010001101001;     //475pi/512
  assign cos2[475]  =  14'b11010011111000;     //475pi/512
  assign sin2[476]  =  14'b11010001110111;     //476pi/512
  assign cos2[476]  =  14'b11010011101001;     //476pi/512
  assign sin2[477]  =  14'b11010010000101;     //477pi/512
  assign cos2[477]  =  14'b11010011011011;     //477pi/512
  assign sin2[478]  =  14'b11010010010011;     //478pi/512
  assign cos2[478]  =  14'b11010011001100;     //478pi/512
  assign sin2[479]  =  14'b11010010100010;     //479pi/512
  assign cos2[479]  =  14'b11010010111110;     //479pi/512
  assign sin2[480]  =  14'b11010010110000;     //480pi/512
  assign cos2[480]  =  14'b11010010110000;     //480pi/512
  assign sin2[481]  =  14'b11010010111110;     //481pi/512
  assign cos2[481]  =  14'b11010010100010;     //481pi/512
  assign sin2[482]  =  14'b11010011001100;     //482pi/512
  assign cos2[482]  =  14'b11010010010011;     //482pi/512
  assign sin2[483]  =  14'b11010011011011;     //483pi/512
  assign cos2[483]  =  14'b11010010000101;     //483pi/512
  assign sin2[484]  =  14'b11010011101001;     //484pi/512
  assign cos2[484]  =  14'b11010001110111;     //484pi/512
  assign sin2[485]  =  14'b11010011111000;     //485pi/512
  assign cos2[485]  =  14'b11010001101001;     //485pi/512
  assign sin2[486]  =  14'b11010100000110;     //486pi/512
  assign cos2[486]  =  14'b11010001011100;     //486pi/512
  assign sin2[487]  =  14'b11010100010101;     //487pi/512
  assign cos2[487]  =  14'b11010001001110;     //487pi/512
  assign sin2[488]  =  14'b11010100100100;     //488pi/512
  assign cos2[488]  =  14'b11010001000000;     //488pi/512
  assign sin2[489]  =  14'b11010100110010;     //489pi/512
  assign cos2[489]  =  14'b11010000110011;     //489pi/512
  assign sin2[490]  =  14'b11010101000001;     //490pi/512
  assign cos2[490]  =  14'b11010000100101;     //490pi/512
  assign sin2[491]  =  14'b11010101010000;     //491pi/512
  assign cos2[491]  =  14'b11010000011000;     //491pi/512
  assign sin2[492]  =  14'b11010101011111;     //492pi/512
  assign cos2[492]  =  14'b11010000001010;     //492pi/512
  assign sin2[493]  =  14'b11010101101110;     //493pi/512
  assign cos2[493]  =  14'b11001111111101;     //493pi/512
  assign sin2[494]  =  14'b11010101111101;     //494pi/512
  assign cos2[494]  =  14'b11001111110000;     //494pi/512
  assign sin2[495]  =  14'b11010110001101;     //495pi/512
  assign cos2[495]  =  14'b11001111100010;     //495pi/512
  assign sin2[496]  =  14'b11010110011100;     //496pi/512
  assign cos2[496]  =  14'b11001111010101;     //496pi/512
  assign sin2[497]  =  14'b11010110101011;     //497pi/512
  assign cos2[497]  =  14'b11001111001000;     //497pi/512
  assign sin2[498]  =  14'b11010110111011;     //498pi/512
  assign cos2[498]  =  14'b11001110111011;     //498pi/512
  assign sin2[499]  =  14'b11010111001010;     //499pi/512
  assign cos2[499]  =  14'b11001110101111;     //499pi/512
  assign sin2[500]  =  14'b11010111011010;     //500pi/512
  assign cos2[500]  =  14'b11001110100010;     //500pi/512
  assign sin2[501]  =  14'b11010111101001;     //501pi/512
  assign cos2[501]  =  14'b11001110010101;     //501pi/512
  assign sin2[502]  =  14'b11010111111001;     //502pi/512
  assign cos2[502]  =  14'b11001110001000;     //502pi/512
  assign sin2[503]  =  14'b11011000001000;     //503pi/512
  assign cos2[503]  =  14'b11001101111100;     //503pi/512
  assign sin2[504]  =  14'b11011000011000;     //504pi/512
  assign cos2[504]  =  14'b11001101101111;     //504pi/512
  assign sin2[505]  =  14'b11011000101000;     //505pi/512
  assign cos2[505]  =  14'b11001101100011;     //505pi/512
  assign sin2[506]  =  14'b11011000111000;     //506pi/512
  assign cos2[506]  =  14'b11001101010111;     //506pi/512
  assign sin2[507]  =  14'b11011001001000;     //507pi/512
  assign cos2[507]  =  14'b11001101001010;     //507pi/512
  assign sin2[508]  =  14'b11011001011000;     //508pi/512
  assign cos2[508]  =  14'b11001100111110;     //508pi/512
  assign sin2[509]  =  14'b11011001101000;     //509pi/512
  assign cos2[509]  =  14'b11001100110010;     //509pi/512
  assign sin2[510]  =  14'b11011001111000;     //510pi/512
  assign cos2[510]  =  14'b11001100100110;     //510pi/512
  assign sin2[511]  =  14'b11011010001000;     //511pi/512
  assign cos2[511]  =  14'b11001100011010;     //511pi/512

endmodule