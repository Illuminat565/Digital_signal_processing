module  M_TWIDLE_12_B_0_10_v  #(parameter SIZE = 10, word_length_tw = 12) (
    input            clk,
    input            en_rd,
    input   [10:0]   rd_ptr_angle,
    input            en_modf,
    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );
reg signed [word_length_tw-1:0]  cos    [511:0];
reg signed [word_length_tw-1:0]  sin    [511:0];
reg signed [word_length_tw-1:0]  m_cos  [511:0];
reg signed [word_length_tw-1:0]  m_sin  [511:0];
reg signed [word_length_tw-1:0]  cos_temp;
reg signed [word_length_tw-1:0]  sin_temp;
reg signed [word_length_tw-1:0]  m_cos_temp;
reg signed [word_length_tw-1:0]  m_sin_temp;
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & ~ en_modf) begin
                  cos_temp           <= cos   [rd_ptr_angle];
                  sin_temp           <= sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & en_modf) begin
                  m_cos_temp           <= m_cos   [rd_ptr_angle];
                  m_sin_temp           <= m_sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(*) begin 
             if (en_modf) begin
                  cos_data           <= m_cos_temp;
                  sin_data           <= m_sin_temp;
             end else begin
                  cos_data           <= cos_temp;
                  sin_data           <= sin_temp;
             end 
        end
initial begin
   sin[0]  =  12'b000000000000;     //0pi/512
   cos[0]  =  12'b010000000000;     //0pi/512
   sin[1]  =  12'b111111111010;     //1pi/512
   cos[1]  =  12'b001111111111;     //1pi/512
   sin[2]  =  12'b111111110011;     //2pi/512
   cos[2]  =  12'b001111111111;     //2pi/512
   sin[3]  =  12'b111111101101;     //3pi/512
   cos[3]  =  12'b001111111111;     //3pi/512
   sin[4]  =  12'b111111100111;     //4pi/512
   cos[4]  =  12'b001111111111;     //4pi/512
   sin[5]  =  12'b111111100001;     //5pi/512
   cos[5]  =  12'b001111111111;     //5pi/512
   sin[6]  =  12'b111111011010;     //6pi/512
   cos[6]  =  12'b001111111111;     //6pi/512
   sin[7]  =  12'b111111010100;     //7pi/512
   cos[7]  =  12'b001111111111;     //7pi/512
   sin[8]  =  12'b111111001110;     //8pi/512
   cos[8]  =  12'b001111111110;     //8pi/512
   sin[9]  =  12'b111111000111;     //9pi/512
   cos[9]  =  12'b001111111110;     //9pi/512
   sin[10]  =  12'b111111000001;     //10pi/512
   cos[10]  =  12'b001111111110;     //10pi/512
   sin[11]  =  12'b111110111011;     //11pi/512
   cos[11]  =  12'b001111111101;     //11pi/512
   sin[12]  =  12'b111110110101;     //12pi/512
   cos[12]  =  12'b001111111101;     //12pi/512
   sin[13]  =  12'b111110101110;     //13pi/512
   cos[13]  =  12'b001111111100;     //13pi/512
   sin[14]  =  12'b111110101000;     //14pi/512
   cos[14]  =  12'b001111111100;     //14pi/512
   sin[15]  =  12'b111110100010;     //15pi/512
   cos[15]  =  12'b001111111011;     //15pi/512
   sin[16]  =  12'b111110011100;     //16pi/512
   cos[16]  =  12'b001111111011;     //16pi/512
   sin[17]  =  12'b111110010101;     //17pi/512
   cos[17]  =  12'b001111111010;     //17pi/512
   sin[18]  =  12'b111110001111;     //18pi/512
   cos[18]  =  12'b001111111001;     //18pi/512
   sin[19]  =  12'b111110001001;     //19pi/512
   cos[19]  =  12'b001111111001;     //19pi/512
   sin[20]  =  12'b111110000011;     //20pi/512
   cos[20]  =  12'b001111111000;     //20pi/512
   sin[21]  =  12'b111101111100;     //21pi/512
   cos[21]  =  12'b001111110111;     //21pi/512
   sin[22]  =  12'b111101110110;     //22pi/512
   cos[22]  =  12'b001111110110;     //22pi/512
   sin[23]  =  12'b111101110000;     //23pi/512
   cos[23]  =  12'b001111110101;     //23pi/512
   sin[24]  =  12'b111101101010;     //24pi/512
   cos[24]  =  12'b001111110100;     //24pi/512
   sin[25]  =  12'b111101100100;     //25pi/512
   cos[25]  =  12'b001111110011;     //25pi/512
   sin[26]  =  12'b111101011101;     //26pi/512
   cos[26]  =  12'b001111110010;     //26pi/512
   sin[27]  =  12'b111101010111;     //27pi/512
   cos[27]  =  12'b001111110001;     //27pi/512
   sin[28]  =  12'b111101010001;     //28pi/512
   cos[28]  =  12'b001111110000;     //28pi/512
   sin[29]  =  12'b111101001011;     //29pi/512
   cos[29]  =  12'b001111101111;     //29pi/512
   sin[30]  =  12'b111101000101;     //30pi/512
   cos[30]  =  12'b001111101110;     //30pi/512
   sin[31]  =  12'b111100111110;     //31pi/512
   cos[31]  =  12'b001111101101;     //31pi/512
   sin[32]  =  12'b111100111000;     //32pi/512
   cos[32]  =  12'b001111101100;     //32pi/512
   sin[33]  =  12'b111100110010;     //33pi/512
   cos[33]  =  12'b001111101011;     //33pi/512
   sin[34]  =  12'b111100101100;     //34pi/512
   cos[34]  =  12'b001111101001;     //34pi/512
   sin[35]  =  12'b111100100110;     //35pi/512
   cos[35]  =  12'b001111101000;     //35pi/512
   sin[36]  =  12'b111100100000;     //36pi/512
   cos[36]  =  12'b001111100111;     //36pi/512
   sin[37]  =  12'b111100011010;     //37pi/512
   cos[37]  =  12'b001111100101;     //37pi/512
   sin[38]  =  12'b111100010011;     //38pi/512
   cos[38]  =  12'b001111100100;     //38pi/512
   sin[39]  =  12'b111100001101;     //39pi/512
   cos[39]  =  12'b001111100010;     //39pi/512
   sin[40]  =  12'b111100000111;     //40pi/512
   cos[40]  =  12'b001111100001;     //40pi/512
   sin[41]  =  12'b111100000001;     //41pi/512
   cos[41]  =  12'b001111011111;     //41pi/512
   sin[42]  =  12'b111011111011;     //42pi/512
   cos[42]  =  12'b001111011110;     //42pi/512
   sin[43]  =  12'b111011110101;     //43pi/512
   cos[43]  =  12'b001111011100;     //43pi/512
   sin[44]  =  12'b111011101111;     //44pi/512
   cos[44]  =  12'b001111011010;     //44pi/512
   sin[45]  =  12'b111011101001;     //45pi/512
   cos[45]  =  12'b001111011001;     //45pi/512
   sin[46]  =  12'b111011100011;     //46pi/512
   cos[46]  =  12'b001111010111;     //46pi/512
   sin[47]  =  12'b111011011101;     //47pi/512
   cos[47]  =  12'b001111010101;     //47pi/512
   sin[48]  =  12'b111011010111;     //48pi/512
   cos[48]  =  12'b001111010011;     //48pi/512
   sin[49]  =  12'b111011010001;     //49pi/512
   cos[49]  =  12'b001111010010;     //49pi/512
   sin[50]  =  12'b111011001011;     //50pi/512
   cos[50]  =  12'b001111010000;     //50pi/512
   sin[51]  =  12'b111011000101;     //51pi/512
   cos[51]  =  12'b001111001110;     //51pi/512
   sin[52]  =  12'b111010111111;     //52pi/512
   cos[52]  =  12'b001111001100;     //52pi/512
   sin[53]  =  12'b111010111001;     //53pi/512
   cos[53]  =  12'b001111001010;     //53pi/512
   sin[54]  =  12'b111010110011;     //54pi/512
   cos[54]  =  12'b001111001000;     //54pi/512
   sin[55]  =  12'b111010101101;     //55pi/512
   cos[55]  =  12'b001111000110;     //55pi/512
   sin[56]  =  12'b111010100111;     //56pi/512
   cos[56]  =  12'b001111000100;     //56pi/512
   sin[57]  =  12'b111010100001;     //57pi/512
   cos[57]  =  12'b001111000010;     //57pi/512
   sin[58]  =  12'b111010011011;     //58pi/512
   cos[58]  =  12'b001110111111;     //58pi/512
   sin[59]  =  12'b111010010101;     //59pi/512
   cos[59]  =  12'b001110111101;     //59pi/512
   sin[60]  =  12'b111010001111;     //60pi/512
   cos[60]  =  12'b001110111011;     //60pi/512
   sin[61]  =  12'b111010001010;     //61pi/512
   cos[61]  =  12'b001110111001;     //61pi/512
   sin[62]  =  12'b111010000100;     //62pi/512
   cos[62]  =  12'b001110110110;     //62pi/512
   sin[63]  =  12'b111001111110;     //63pi/512
   cos[63]  =  12'b001110110100;     //63pi/512
   sin[64]  =  12'b111001111000;     //64pi/512
   cos[64]  =  12'b001110110010;     //64pi/512
   sin[65]  =  12'b111001110010;     //65pi/512
   cos[65]  =  12'b001110101111;     //65pi/512
   sin[66]  =  12'b111001101101;     //66pi/512
   cos[66]  =  12'b001110101101;     //66pi/512
   sin[67]  =  12'b111001100111;     //67pi/512
   cos[67]  =  12'b001110101010;     //67pi/512
   sin[68]  =  12'b111001100001;     //68pi/512
   cos[68]  =  12'b001110101000;     //68pi/512
   sin[69]  =  12'b111001011011;     //69pi/512
   cos[69]  =  12'b001110100101;     //69pi/512
   sin[70]  =  12'b111001010110;     //70pi/512
   cos[70]  =  12'b001110100010;     //70pi/512
   sin[71]  =  12'b111001010000;     //71pi/512
   cos[71]  =  12'b001110100000;     //71pi/512
   sin[72]  =  12'b111001001010;     //72pi/512
   cos[72]  =  12'b001110011101;     //72pi/512
   sin[73]  =  12'b111001000101;     //73pi/512
   cos[73]  =  12'b001110011010;     //73pi/512
   sin[74]  =  12'b111000111111;     //74pi/512
   cos[74]  =  12'b001110011000;     //74pi/512
   sin[75]  =  12'b111000111001;     //75pi/512
   cos[75]  =  12'b001110010101;     //75pi/512
   sin[76]  =  12'b111000110100;     //76pi/512
   cos[76]  =  12'b001110010010;     //76pi/512
   sin[77]  =  12'b111000101110;     //77pi/512
   cos[77]  =  12'b001110001111;     //77pi/512
   sin[78]  =  12'b111000101000;     //78pi/512
   cos[78]  =  12'b001110001100;     //78pi/512
   sin[79]  =  12'b111000100011;     //79pi/512
   cos[79]  =  12'b001110001010;     //79pi/512
   sin[80]  =  12'b111000011101;     //80pi/512
   cos[80]  =  12'b001110000111;     //80pi/512
   sin[81]  =  12'b111000011000;     //81pi/512
   cos[81]  =  12'b001110000100;     //81pi/512
   sin[82]  =  12'b111000010010;     //82pi/512
   cos[82]  =  12'b001110000001;     //82pi/512
   sin[83]  =  12'b111000001101;     //83pi/512
   cos[83]  =  12'b001101111110;     //83pi/512
   sin[84]  =  12'b111000000111;     //84pi/512
   cos[84]  =  12'b001101111010;     //84pi/512
   sin[85]  =  12'b111000000010;     //85pi/512
   cos[85]  =  12'b001101110111;     //85pi/512
   sin[86]  =  12'b110111111100;     //86pi/512
   cos[86]  =  12'b001101110100;     //86pi/512
   sin[87]  =  12'b110111110111;     //87pi/512
   cos[87]  =  12'b001101110001;     //87pi/512
   sin[88]  =  12'b110111110010;     //88pi/512
   cos[88]  =  12'b001101101110;     //88pi/512
   sin[89]  =  12'b110111101100;     //89pi/512
   cos[89]  =  12'b001101101011;     //89pi/512
   sin[90]  =  12'b110111100111;     //90pi/512
   cos[90]  =  12'b001101100111;     //90pi/512
   sin[91]  =  12'b110111100001;     //91pi/512
   cos[91]  =  12'b001101100100;     //91pi/512
   sin[92]  =  12'b110111011100;     //92pi/512
   cos[92]  =  12'b001101100001;     //92pi/512
   sin[93]  =  12'b110111010111;     //93pi/512
   cos[93]  =  12'b001101011101;     //93pi/512
   sin[94]  =  12'b110111010010;     //94pi/512
   cos[94]  =  12'b001101011010;     //94pi/512
   sin[95]  =  12'b110111001100;     //95pi/512
   cos[95]  =  12'b001101010110;     //95pi/512
   sin[96]  =  12'b110111000111;     //96pi/512
   cos[96]  =  12'b001101010011;     //96pi/512
   sin[97]  =  12'b110111000010;     //97pi/512
   cos[97]  =  12'b001101001111;     //97pi/512
   sin[98]  =  12'b110110111101;     //98pi/512
   cos[98]  =  12'b001101001100;     //98pi/512
   sin[99]  =  12'b110110111000;     //99pi/512
   cos[99]  =  12'b001101001000;     //99pi/512
   sin[100]  =  12'b110110110010;     //100pi/512
   cos[100]  =  12'b001101000101;     //100pi/512
   sin[101]  =  12'b110110101101;     //101pi/512
   cos[101]  =  12'b001101000001;     //101pi/512
   sin[102]  =  12'b110110101000;     //102pi/512
   cos[102]  =  12'b001100111101;     //102pi/512
   sin[103]  =  12'b110110100011;     //103pi/512
   cos[103]  =  12'b001100111010;     //103pi/512
   sin[104]  =  12'b110110011110;     //104pi/512
   cos[104]  =  12'b001100110110;     //104pi/512
   sin[105]  =  12'b110110011001;     //105pi/512
   cos[105]  =  12'b001100110010;     //105pi/512
   sin[106]  =  12'b110110010100;     //106pi/512
   cos[106]  =  12'b001100101110;     //106pi/512
   sin[107]  =  12'b110110001111;     //107pi/512
   cos[107]  =  12'b001100101011;     //107pi/512
   sin[108]  =  12'b110110001010;     //108pi/512
   cos[108]  =  12'b001100100111;     //108pi/512
   sin[109]  =  12'b110110000101;     //109pi/512
   cos[109]  =  12'b001100100011;     //109pi/512
   sin[110]  =  12'b110110000000;     //110pi/512
   cos[110]  =  12'b001100011111;     //110pi/512
   sin[111]  =  12'b110101111011;     //111pi/512
   cos[111]  =  12'b001100011011;     //111pi/512
   sin[112]  =  12'b110101110110;     //112pi/512
   cos[112]  =  12'b001100010111;     //112pi/512
   sin[113]  =  12'b110101110010;     //113pi/512
   cos[113]  =  12'b001100010011;     //113pi/512
   sin[114]  =  12'b110101101101;     //114pi/512
   cos[114]  =  12'b001100001111;     //114pi/512
   sin[115]  =  12'b110101101000;     //115pi/512
   cos[115]  =  12'b001100001011;     //115pi/512
   sin[116]  =  12'b110101100011;     //116pi/512
   cos[116]  =  12'b001100000111;     //116pi/512
   sin[117]  =  12'b110101011110;     //117pi/512
   cos[117]  =  12'b001100000011;     //117pi/512
   sin[118]  =  12'b110101011010;     //118pi/512
   cos[118]  =  12'b001011111111;     //118pi/512
   sin[119]  =  12'b110101010101;     //119pi/512
   cos[119]  =  12'b001011111010;     //119pi/512
   sin[120]  =  12'b110101010000;     //120pi/512
   cos[120]  =  12'b001011110110;     //120pi/512
   sin[121]  =  12'b110101001100;     //121pi/512
   cos[121]  =  12'b001011110010;     //121pi/512
   sin[122]  =  12'b110101000111;     //122pi/512
   cos[122]  =  12'b001011101110;     //122pi/512
   sin[123]  =  12'b110101000010;     //123pi/512
   cos[123]  =  12'b001011101001;     //123pi/512
   sin[124]  =  12'b110100111110;     //124pi/512
   cos[124]  =  12'b001011100101;     //124pi/512
   sin[125]  =  12'b110100111001;     //125pi/512
   cos[125]  =  12'b001011100001;     //125pi/512
   sin[126]  =  12'b110100110101;     //126pi/512
   cos[126]  =  12'b001011011100;     //126pi/512
   sin[127]  =  12'b110100110000;     //127pi/512
   cos[127]  =  12'b001011011000;     //127pi/512
   sin[128]  =  12'b110100101100;     //128pi/512
   cos[128]  =  12'b001011010100;     //128pi/512
   sin[129]  =  12'b110100100111;     //129pi/512
   cos[129]  =  12'b001011001111;     //129pi/512
   sin[130]  =  12'b110100100011;     //130pi/512
   cos[130]  =  12'b001011001011;     //130pi/512
   sin[131]  =  12'b110100011111;     //131pi/512
   cos[131]  =  12'b001011000110;     //131pi/512
   sin[132]  =  12'b110100011010;     //132pi/512
   cos[132]  =  12'b001011000010;     //132pi/512
   sin[133]  =  12'b110100010110;     //133pi/512
   cos[133]  =  12'b001010111101;     //133pi/512
   sin[134]  =  12'b110100010010;     //134pi/512
   cos[134]  =  12'b001010111000;     //134pi/512
   sin[135]  =  12'b110100001101;     //135pi/512
   cos[135]  =  12'b001010110100;     //135pi/512
   sin[136]  =  12'b110100001001;     //136pi/512
   cos[136]  =  12'b001010101111;     //136pi/512
   sin[137]  =  12'b110100000101;     //137pi/512
   cos[137]  =  12'b001010101011;     //137pi/512
   sin[138]  =  12'b110100000001;     //138pi/512
   cos[138]  =  12'b001010100110;     //138pi/512
   sin[139]  =  12'b110011111101;     //139pi/512
   cos[139]  =  12'b001010100001;     //139pi/512
   sin[140]  =  12'b110011111001;     //140pi/512
   cos[140]  =  12'b001010011100;     //140pi/512
   sin[141]  =  12'b110011110101;     //141pi/512
   cos[141]  =  12'b001010011000;     //141pi/512
   sin[142]  =  12'b110011110000;     //142pi/512
   cos[142]  =  12'b001010010011;     //142pi/512
   sin[143]  =  12'b110011101100;     //143pi/512
   cos[143]  =  12'b001010001110;     //143pi/512
   sin[144]  =  12'b110011101000;     //144pi/512
   cos[144]  =  12'b001010001001;     //144pi/512
   sin[145]  =  12'b110011100100;     //145pi/512
   cos[145]  =  12'b001010000100;     //145pi/512
   sin[146]  =  12'b110011100001;     //146pi/512
   cos[146]  =  12'b001001111111;     //146pi/512
   sin[147]  =  12'b110011011101;     //147pi/512
   cos[147]  =  12'b001001111010;     //147pi/512
   sin[148]  =  12'b110011011001;     //148pi/512
   cos[148]  =  12'b001001110101;     //148pi/512
   sin[149]  =  12'b110011010101;     //149pi/512
   cos[149]  =  12'b001001110001;     //149pi/512
   sin[150]  =  12'b110011010001;     //150pi/512
   cos[150]  =  12'b001001101100;     //150pi/512
   sin[151]  =  12'b110011001101;     //151pi/512
   cos[151]  =  12'b001001100111;     //151pi/512
   sin[152]  =  12'b110011001010;     //152pi/512
   cos[152]  =  12'b001001100001;     //152pi/512
   sin[153]  =  12'b110011000110;     //153pi/512
   cos[153]  =  12'b001001011100;     //153pi/512
   sin[154]  =  12'b110011000010;     //154pi/512
   cos[154]  =  12'b001001010111;     //154pi/512
   sin[155]  =  12'b110010111110;     //155pi/512
   cos[155]  =  12'b001001010010;     //155pi/512
   sin[156]  =  12'b110010111011;     //156pi/512
   cos[156]  =  12'b001001001101;     //156pi/512
   sin[157]  =  12'b110010110111;     //157pi/512
   cos[157]  =  12'b001001001000;     //157pi/512
   sin[158]  =  12'b110010110100;     //158pi/512
   cos[158]  =  12'b001001000011;     //158pi/512
   sin[159]  =  12'b110010110000;     //159pi/512
   cos[159]  =  12'b001000111110;     //159pi/512
   sin[160]  =  12'b110010101101;     //160pi/512
   cos[160]  =  12'b001000111000;     //160pi/512
   sin[161]  =  12'b110010101001;     //161pi/512
   cos[161]  =  12'b001000110011;     //161pi/512
   sin[162]  =  12'b110010100110;     //162pi/512
   cos[162]  =  12'b001000101110;     //162pi/512
   sin[163]  =  12'b110010100010;     //163pi/512
   cos[163]  =  12'b001000101001;     //163pi/512
   sin[164]  =  12'b110010011111;     //164pi/512
   cos[164]  =  12'b001000100011;     //164pi/512
   sin[165]  =  12'b110010011100;     //165pi/512
   cos[165]  =  12'b001000011110;     //165pi/512
   sin[166]  =  12'b110010011000;     //166pi/512
   cos[166]  =  12'b001000011001;     //166pi/512
   sin[167]  =  12'b110010010101;     //167pi/512
   cos[167]  =  12'b001000010011;     //167pi/512
   sin[168]  =  12'b110010010010;     //168pi/512
   cos[168]  =  12'b001000001110;     //168pi/512
   sin[169]  =  12'b110010001110;     //169pi/512
   cos[169]  =  12'b001000001001;     //169pi/512
   sin[170]  =  12'b110010001011;     //170pi/512
   cos[170]  =  12'b001000000011;     //170pi/512
   sin[171]  =  12'b110010001000;     //171pi/512
   cos[171]  =  12'b000111111110;     //171pi/512
   sin[172]  =  12'b110010000101;     //172pi/512
   cos[172]  =  12'b000111111000;     //172pi/512
   sin[173]  =  12'b110010000010;     //173pi/512
   cos[173]  =  12'b000111110011;     //173pi/512
   sin[174]  =  12'b110001111111;     //174pi/512
   cos[174]  =  12'b000111101101;     //174pi/512
   sin[175]  =  12'b110001111100;     //175pi/512
   cos[175]  =  12'b000111101000;     //175pi/512
   sin[176]  =  12'b110001111001;     //176pi/512
   cos[176]  =  12'b000111100010;     //176pi/512
   sin[177]  =  12'b110001110110;     //177pi/512
   cos[177]  =  12'b000111011101;     //177pi/512
   sin[178]  =  12'b110001110011;     //178pi/512
   cos[178]  =  12'b000111010111;     //178pi/512
   sin[179]  =  12'b110001110000;     //179pi/512
   cos[179]  =  12'b000111010010;     //179pi/512
   sin[180]  =  12'b110001101101;     //180pi/512
   cos[180]  =  12'b000111001100;     //180pi/512
   sin[181]  =  12'b110001101011;     //181pi/512
   cos[181]  =  12'b000111000110;     //181pi/512
   sin[182]  =  12'b110001101000;     //182pi/512
   cos[182]  =  12'b000111000001;     //182pi/512
   sin[183]  =  12'b110001100101;     //183pi/512
   cos[183]  =  12'b000110111011;     //183pi/512
   sin[184]  =  12'b110001100010;     //184pi/512
   cos[184]  =  12'b000110110101;     //184pi/512
   sin[185]  =  12'b110001100000;     //185pi/512
   cos[185]  =  12'b000110110000;     //185pi/512
   sin[186]  =  12'b110001011101;     //186pi/512
   cos[186]  =  12'b000110101010;     //186pi/512
   sin[187]  =  12'b110001011010;     //187pi/512
   cos[187]  =  12'b000110100100;     //187pi/512
   sin[188]  =  12'b110001011000;     //188pi/512
   cos[188]  =  12'b000110011110;     //188pi/512
   sin[189]  =  12'b110001010101;     //189pi/512
   cos[189]  =  12'b000110011001;     //189pi/512
   sin[190]  =  12'b110001010011;     //190pi/512
   cos[190]  =  12'b000110010011;     //190pi/512
   sin[191]  =  12'b110001010000;     //191pi/512
   cos[191]  =  12'b000110001101;     //191pi/512
   sin[192]  =  12'b110001001110;     //192pi/512
   cos[192]  =  12'b000110000111;     //192pi/512
   sin[193]  =  12'b110001001100;     //193pi/512
   cos[193]  =  12'b000110000010;     //193pi/512
   sin[194]  =  12'b110001001001;     //194pi/512
   cos[194]  =  12'b000101111100;     //194pi/512
   sin[195]  =  12'b110001000111;     //195pi/512
   cos[195]  =  12'b000101110110;     //195pi/512
   sin[196]  =  12'b110001000101;     //196pi/512
   cos[196]  =  12'b000101110000;     //196pi/512
   sin[197]  =  12'b110001000010;     //197pi/512
   cos[197]  =  12'b000101101010;     //197pi/512
   sin[198]  =  12'b110001000000;     //198pi/512
   cos[198]  =  12'b000101100100;     //198pi/512
   sin[199]  =  12'b110000111110;     //199pi/512
   cos[199]  =  12'b000101011110;     //199pi/512
   sin[200]  =  12'b110000111100;     //200pi/512
   cos[200]  =  12'b000101011000;     //200pi/512
   sin[201]  =  12'b110000111010;     //201pi/512
   cos[201]  =  12'b000101010011;     //201pi/512
   sin[202]  =  12'b110000111000;     //202pi/512
   cos[202]  =  12'b000101001101;     //202pi/512
   sin[203]  =  12'b110000110110;     //203pi/512
   cos[203]  =  12'b000101000111;     //203pi/512
   sin[204]  =  12'b110000110100;     //204pi/512
   cos[204]  =  12'b000101000001;     //204pi/512
   sin[205]  =  12'b110000110010;     //205pi/512
   cos[205]  =  12'b000100111011;     //205pi/512
   sin[206]  =  12'b110000110000;     //206pi/512
   cos[206]  =  12'b000100110101;     //206pi/512
   sin[207]  =  12'b110000101110;     //207pi/512
   cos[207]  =  12'b000100101111;     //207pi/512
   sin[208]  =  12'b110000101100;     //208pi/512
   cos[208]  =  12'b000100101001;     //208pi/512
   sin[209]  =  12'b110000101010;     //209pi/512
   cos[209]  =  12'b000100100011;     //209pi/512
   sin[210]  =  12'b110000101001;     //210pi/512
   cos[210]  =  12'b000100011101;     //210pi/512
   sin[211]  =  12'b110000100111;     //211pi/512
   cos[211]  =  12'b000100010111;     //211pi/512
   sin[212]  =  12'b110000100101;     //212pi/512
   cos[212]  =  12'b000100010001;     //212pi/512
   sin[213]  =  12'b110000100011;     //213pi/512
   cos[213]  =  12'b000100001011;     //213pi/512
   sin[214]  =  12'b110000100010;     //214pi/512
   cos[214]  =  12'b000100000100;     //214pi/512
   sin[215]  =  12'b110000100000;     //215pi/512
   cos[215]  =  12'b000011111110;     //215pi/512
   sin[216]  =  12'b110000011111;     //216pi/512
   cos[216]  =  12'b000011111000;     //216pi/512
   sin[217]  =  12'b110000011101;     //217pi/512
   cos[217]  =  12'b000011110010;     //217pi/512
   sin[218]  =  12'b110000011100;     //218pi/512
   cos[218]  =  12'b000011101100;     //218pi/512
   sin[219]  =  12'b110000011010;     //219pi/512
   cos[219]  =  12'b000011100110;     //219pi/512
   sin[220]  =  12'b110000011001;     //220pi/512
   cos[220]  =  12'b000011100000;     //220pi/512
   sin[221]  =  12'b110000011000;     //221pi/512
   cos[221]  =  12'b000011011010;     //221pi/512
   sin[222]  =  12'b110000010110;     //222pi/512
   cos[222]  =  12'b000011010100;     //222pi/512
   sin[223]  =  12'b110000010101;     //223pi/512
   cos[223]  =  12'b000011001101;     //223pi/512
   sin[224]  =  12'b110000010100;     //224pi/512
   cos[224]  =  12'b000011000111;     //224pi/512
   sin[225]  =  12'b110000010010;     //225pi/512
   cos[225]  =  12'b000011000001;     //225pi/512
   sin[226]  =  12'b110000010001;     //226pi/512
   cos[226]  =  12'b000010111011;     //226pi/512
   sin[227]  =  12'b110000010000;     //227pi/512
   cos[227]  =  12'b000010110101;     //227pi/512
   sin[228]  =  12'b110000001111;     //228pi/512
   cos[228]  =  12'b000010101111;     //228pi/512
   sin[229]  =  12'b110000001110;     //229pi/512
   cos[229]  =  12'b000010101000;     //229pi/512
   sin[230]  =  12'b110000001101;     //230pi/512
   cos[230]  =  12'b000010100010;     //230pi/512
   sin[231]  =  12'b110000001100;     //231pi/512
   cos[231]  =  12'b000010011100;     //231pi/512
   sin[232]  =  12'b110000001011;     //232pi/512
   cos[232]  =  12'b000010010110;     //232pi/512
   sin[233]  =  12'b110000001010;     //233pi/512
   cos[233]  =  12'b000010010000;     //233pi/512
   sin[234]  =  12'b110000001001;     //234pi/512
   cos[234]  =  12'b000010001001;     //234pi/512
   sin[235]  =  12'b110000001000;     //235pi/512
   cos[235]  =  12'b000010000011;     //235pi/512
   sin[236]  =  12'b110000001000;     //236pi/512
   cos[236]  =  12'b000001111101;     //236pi/512
   sin[237]  =  12'b110000000111;     //237pi/512
   cos[237]  =  12'b000001110111;     //237pi/512
   sin[238]  =  12'b110000000110;     //238pi/512
   cos[238]  =  12'b000001110000;     //238pi/512
   sin[239]  =  12'b110000000110;     //239pi/512
   cos[239]  =  12'b000001101010;     //239pi/512
   sin[240]  =  12'b110000000101;     //240pi/512
   cos[240]  =  12'b000001100100;     //240pi/512
   sin[241]  =  12'b110000000100;     //241pi/512
   cos[241]  =  12'b000001011110;     //241pi/512
   sin[242]  =  12'b110000000100;     //242pi/512
   cos[242]  =  12'b000001010111;     //242pi/512
   sin[243]  =  12'b110000000011;     //243pi/512
   cos[243]  =  12'b000001010001;     //243pi/512
   sin[244]  =  12'b110000000011;     //244pi/512
   cos[244]  =  12'b000001001011;     //244pi/512
   sin[245]  =  12'b110000000010;     //245pi/512
   cos[245]  =  12'b000001000101;     //245pi/512
   sin[246]  =  12'b110000000010;     //246pi/512
   cos[246]  =  12'b000000111110;     //246pi/512
   sin[247]  =  12'b110000000010;     //247pi/512
   cos[247]  =  12'b000000111000;     //247pi/512
   sin[248]  =  12'b110000000001;     //248pi/512
   cos[248]  =  12'b000000110010;     //248pi/512
   sin[249]  =  12'b110000000001;     //249pi/512
   cos[249]  =  12'b000000101011;     //249pi/512
   sin[250]  =  12'b110000000001;     //250pi/512
   cos[250]  =  12'b000000100101;     //250pi/512
   sin[251]  =  12'b110000000000;     //251pi/512
   cos[251]  =  12'b000000011111;     //251pi/512
   sin[252]  =  12'b110000000000;     //252pi/512
   cos[252]  =  12'b000000011001;     //252pi/512
   sin[253]  =  12'b110000000000;     //253pi/512
   cos[253]  =  12'b000000010010;     //253pi/512
   sin[254]  =  12'b110000000000;     //254pi/512
   cos[254]  =  12'b000000001100;     //254pi/512
   sin[255]  =  12'b110000000000;     //255pi/512
   cos[255]  =  12'b000000000110;     //255pi/512
   sin[256]  =  12'b110000000000;     //256pi/512
   cos[256]  =  12'b000000000000;     //256pi/512
   sin[257]  =  12'b110000000000;     //257pi/512
   cos[257]  =  12'b111111111010;     //257pi/512
   sin[258]  =  12'b110000000000;     //258pi/512
   cos[258]  =  12'b111111110011;     //258pi/512
   sin[259]  =  12'b110000000000;     //259pi/512
   cos[259]  =  12'b111111101101;     //259pi/512
   sin[260]  =  12'b110000000000;     //260pi/512
   cos[260]  =  12'b111111100111;     //260pi/512
   sin[261]  =  12'b110000000000;     //261pi/512
   cos[261]  =  12'b111111100001;     //261pi/512
   sin[262]  =  12'b110000000001;     //262pi/512
   cos[262]  =  12'b111111011010;     //262pi/512
   sin[263]  =  12'b110000000001;     //263pi/512
   cos[263]  =  12'b111111010100;     //263pi/512
   sin[264]  =  12'b110000000001;     //264pi/512
   cos[264]  =  12'b111111001110;     //264pi/512
   sin[265]  =  12'b110000000010;     //265pi/512
   cos[265]  =  12'b111111000111;     //265pi/512
   sin[266]  =  12'b110000000010;     //266pi/512
   cos[266]  =  12'b111111000001;     //266pi/512
   sin[267]  =  12'b110000000010;     //267pi/512
   cos[267]  =  12'b111110111011;     //267pi/512
   sin[268]  =  12'b110000000011;     //268pi/512
   cos[268]  =  12'b111110110101;     //268pi/512
   sin[269]  =  12'b110000000011;     //269pi/512
   cos[269]  =  12'b111110101110;     //269pi/512
   sin[270]  =  12'b110000000100;     //270pi/512
   cos[270]  =  12'b111110101000;     //270pi/512
   sin[271]  =  12'b110000000100;     //271pi/512
   cos[271]  =  12'b111110100010;     //271pi/512
   sin[272]  =  12'b110000000101;     //272pi/512
   cos[272]  =  12'b111110011100;     //272pi/512
   sin[273]  =  12'b110000000110;     //273pi/512
   cos[273]  =  12'b111110010101;     //273pi/512
   sin[274]  =  12'b110000000110;     //274pi/512
   cos[274]  =  12'b111110001111;     //274pi/512
   sin[275]  =  12'b110000000111;     //275pi/512
   cos[275]  =  12'b111110001001;     //275pi/512
   sin[276]  =  12'b110000001000;     //276pi/512
   cos[276]  =  12'b111110000011;     //276pi/512
   sin[277]  =  12'b110000001000;     //277pi/512
   cos[277]  =  12'b111101111100;     //277pi/512
   sin[278]  =  12'b110000001001;     //278pi/512
   cos[278]  =  12'b111101110110;     //278pi/512
   sin[279]  =  12'b110000001010;     //279pi/512
   cos[279]  =  12'b111101110000;     //279pi/512
   sin[280]  =  12'b110000001011;     //280pi/512
   cos[280]  =  12'b111101101010;     //280pi/512
   sin[281]  =  12'b110000001100;     //281pi/512
   cos[281]  =  12'b111101100100;     //281pi/512
   sin[282]  =  12'b110000001101;     //282pi/512
   cos[282]  =  12'b111101011101;     //282pi/512
   sin[283]  =  12'b110000001110;     //283pi/512
   cos[283]  =  12'b111101010111;     //283pi/512
   sin[284]  =  12'b110000001111;     //284pi/512
   cos[284]  =  12'b111101010001;     //284pi/512
   sin[285]  =  12'b110000010000;     //285pi/512
   cos[285]  =  12'b111101001011;     //285pi/512
   sin[286]  =  12'b110000010001;     //286pi/512
   cos[286]  =  12'b111101000101;     //286pi/512
   sin[287]  =  12'b110000010010;     //287pi/512
   cos[287]  =  12'b111100111110;     //287pi/512
   sin[288]  =  12'b110000010100;     //288pi/512
   cos[288]  =  12'b111100111000;     //288pi/512
   sin[289]  =  12'b110000010101;     //289pi/512
   cos[289]  =  12'b111100110010;     //289pi/512
   sin[290]  =  12'b110000010110;     //290pi/512
   cos[290]  =  12'b111100101100;     //290pi/512
   sin[291]  =  12'b110000011000;     //291pi/512
   cos[291]  =  12'b111100100110;     //291pi/512
   sin[292]  =  12'b110000011001;     //292pi/512
   cos[292]  =  12'b111100100000;     //292pi/512
   sin[293]  =  12'b110000011010;     //293pi/512
   cos[293]  =  12'b111100011010;     //293pi/512
   sin[294]  =  12'b110000011100;     //294pi/512
   cos[294]  =  12'b111100010011;     //294pi/512
   sin[295]  =  12'b110000011101;     //295pi/512
   cos[295]  =  12'b111100001101;     //295pi/512
   sin[296]  =  12'b110000011111;     //296pi/512
   cos[296]  =  12'b111100000111;     //296pi/512
   sin[297]  =  12'b110000100000;     //297pi/512
   cos[297]  =  12'b111100000001;     //297pi/512
   sin[298]  =  12'b110000100010;     //298pi/512
   cos[298]  =  12'b111011111011;     //298pi/512
   sin[299]  =  12'b110000100011;     //299pi/512
   cos[299]  =  12'b111011110101;     //299pi/512
   sin[300]  =  12'b110000100101;     //300pi/512
   cos[300]  =  12'b111011101111;     //300pi/512
   sin[301]  =  12'b110000100111;     //301pi/512
   cos[301]  =  12'b111011101001;     //301pi/512
   sin[302]  =  12'b110000101001;     //302pi/512
   cos[302]  =  12'b111011100011;     //302pi/512
   sin[303]  =  12'b110000101010;     //303pi/512
   cos[303]  =  12'b111011011101;     //303pi/512
   sin[304]  =  12'b110000101100;     //304pi/512
   cos[304]  =  12'b111011010111;     //304pi/512
   sin[305]  =  12'b110000101110;     //305pi/512
   cos[305]  =  12'b111011010001;     //305pi/512
   sin[306]  =  12'b110000110000;     //306pi/512
   cos[306]  =  12'b111011001011;     //306pi/512
   sin[307]  =  12'b110000110010;     //307pi/512
   cos[307]  =  12'b111011000101;     //307pi/512
   sin[308]  =  12'b110000110100;     //308pi/512
   cos[308]  =  12'b111010111111;     //308pi/512
   sin[309]  =  12'b110000110110;     //309pi/512
   cos[309]  =  12'b111010111001;     //309pi/512
   sin[310]  =  12'b110000111000;     //310pi/512
   cos[310]  =  12'b111010110011;     //310pi/512
   sin[311]  =  12'b110000111010;     //311pi/512
   cos[311]  =  12'b111010101101;     //311pi/512
   sin[312]  =  12'b110000111100;     //312pi/512
   cos[312]  =  12'b111010100111;     //312pi/512
   sin[313]  =  12'b110000111110;     //313pi/512
   cos[313]  =  12'b111010100001;     //313pi/512
   sin[314]  =  12'b110001000000;     //314pi/512
   cos[314]  =  12'b111010011011;     //314pi/512
   sin[315]  =  12'b110001000010;     //315pi/512
   cos[315]  =  12'b111010010101;     //315pi/512
   sin[316]  =  12'b110001000101;     //316pi/512
   cos[316]  =  12'b111010001111;     //316pi/512
   sin[317]  =  12'b110001000111;     //317pi/512
   cos[317]  =  12'b111010001010;     //317pi/512
   sin[318]  =  12'b110001001001;     //318pi/512
   cos[318]  =  12'b111010000100;     //318pi/512
   sin[319]  =  12'b110001001100;     //319pi/512
   cos[319]  =  12'b111001111110;     //319pi/512
   sin[320]  =  12'b110001001110;     //320pi/512
   cos[320]  =  12'b111001111000;     //320pi/512
   sin[321]  =  12'b110001010000;     //321pi/512
   cos[321]  =  12'b111001110010;     //321pi/512
   sin[322]  =  12'b110001010011;     //322pi/512
   cos[322]  =  12'b111001101101;     //322pi/512
   sin[323]  =  12'b110001010101;     //323pi/512
   cos[323]  =  12'b111001100111;     //323pi/512
   sin[324]  =  12'b110001011000;     //324pi/512
   cos[324]  =  12'b111001100001;     //324pi/512
   sin[325]  =  12'b110001011010;     //325pi/512
   cos[325]  =  12'b111001011011;     //325pi/512
   sin[326]  =  12'b110001011101;     //326pi/512
   cos[326]  =  12'b111001010110;     //326pi/512
   sin[327]  =  12'b110001100000;     //327pi/512
   cos[327]  =  12'b111001010000;     //327pi/512
   sin[328]  =  12'b110001100010;     //328pi/512
   cos[328]  =  12'b111001001010;     //328pi/512
   sin[329]  =  12'b110001100101;     //329pi/512
   cos[329]  =  12'b111001000101;     //329pi/512
   sin[330]  =  12'b110001101000;     //330pi/512
   cos[330]  =  12'b111000111111;     //330pi/512
   sin[331]  =  12'b110001101011;     //331pi/512
   cos[331]  =  12'b111000111001;     //331pi/512
   sin[332]  =  12'b110001101101;     //332pi/512
   cos[332]  =  12'b111000110100;     //332pi/512
   sin[333]  =  12'b110001110000;     //333pi/512
   cos[333]  =  12'b111000101110;     //333pi/512
   sin[334]  =  12'b110001110011;     //334pi/512
   cos[334]  =  12'b111000101000;     //334pi/512
   sin[335]  =  12'b110001110110;     //335pi/512
   cos[335]  =  12'b111000100011;     //335pi/512
   sin[336]  =  12'b110001111001;     //336pi/512
   cos[336]  =  12'b111000011101;     //336pi/512
   sin[337]  =  12'b110001111100;     //337pi/512
   cos[337]  =  12'b111000011000;     //337pi/512
   sin[338]  =  12'b110001111111;     //338pi/512
   cos[338]  =  12'b111000010010;     //338pi/512
   sin[339]  =  12'b110010000010;     //339pi/512
   cos[339]  =  12'b111000001101;     //339pi/512
   sin[340]  =  12'b110010000101;     //340pi/512
   cos[340]  =  12'b111000000111;     //340pi/512
   sin[341]  =  12'b110010001000;     //341pi/512
   cos[341]  =  12'b111000000010;     //341pi/512
   sin[342]  =  12'b110010001011;     //342pi/512
   cos[342]  =  12'b110111111100;     //342pi/512
   sin[343]  =  12'b110010001110;     //343pi/512
   cos[343]  =  12'b110111110111;     //343pi/512
   sin[344]  =  12'b110010010010;     //344pi/512
   cos[344]  =  12'b110111110010;     //344pi/512
   sin[345]  =  12'b110010010101;     //345pi/512
   cos[345]  =  12'b110111101100;     //345pi/512
   sin[346]  =  12'b110010011000;     //346pi/512
   cos[346]  =  12'b110111100111;     //346pi/512
   sin[347]  =  12'b110010011100;     //347pi/512
   cos[347]  =  12'b110111100001;     //347pi/512
   sin[348]  =  12'b110010011111;     //348pi/512
   cos[348]  =  12'b110111011100;     //348pi/512
   sin[349]  =  12'b110010100010;     //349pi/512
   cos[349]  =  12'b110111010111;     //349pi/512
   sin[350]  =  12'b110010100110;     //350pi/512
   cos[350]  =  12'b110111010010;     //350pi/512
   sin[351]  =  12'b110010101001;     //351pi/512
   cos[351]  =  12'b110111001100;     //351pi/512
   sin[352]  =  12'b110010101101;     //352pi/512
   cos[352]  =  12'b110111000111;     //352pi/512
   sin[353]  =  12'b110010110000;     //353pi/512
   cos[353]  =  12'b110111000010;     //353pi/512
   sin[354]  =  12'b110010110100;     //354pi/512
   cos[354]  =  12'b110110111101;     //354pi/512
   sin[355]  =  12'b110010110111;     //355pi/512
   cos[355]  =  12'b110110111000;     //355pi/512
   sin[356]  =  12'b110010111011;     //356pi/512
   cos[356]  =  12'b110110110010;     //356pi/512
   sin[357]  =  12'b110010111110;     //357pi/512
   cos[357]  =  12'b110110101101;     //357pi/512
   sin[358]  =  12'b110011000010;     //358pi/512
   cos[358]  =  12'b110110101000;     //358pi/512
   sin[359]  =  12'b110011000110;     //359pi/512
   cos[359]  =  12'b110110100011;     //359pi/512
   sin[360]  =  12'b110011001010;     //360pi/512
   cos[360]  =  12'b110110011110;     //360pi/512
   sin[361]  =  12'b110011001101;     //361pi/512
   cos[361]  =  12'b110110011001;     //361pi/512
   sin[362]  =  12'b110011010001;     //362pi/512
   cos[362]  =  12'b110110010100;     //362pi/512
   sin[363]  =  12'b110011010101;     //363pi/512
   cos[363]  =  12'b110110001111;     //363pi/512
   sin[364]  =  12'b110011011001;     //364pi/512
   cos[364]  =  12'b110110001010;     //364pi/512
   sin[365]  =  12'b110011011101;     //365pi/512
   cos[365]  =  12'b110110000101;     //365pi/512
   sin[366]  =  12'b110011100001;     //366pi/512
   cos[366]  =  12'b110110000000;     //366pi/512
   sin[367]  =  12'b110011100100;     //367pi/512
   cos[367]  =  12'b110101111011;     //367pi/512
   sin[368]  =  12'b110011101000;     //368pi/512
   cos[368]  =  12'b110101110110;     //368pi/512
   sin[369]  =  12'b110011101100;     //369pi/512
   cos[369]  =  12'b110101110010;     //369pi/512
   sin[370]  =  12'b110011110000;     //370pi/512
   cos[370]  =  12'b110101101101;     //370pi/512
   sin[371]  =  12'b110011110101;     //371pi/512
   cos[371]  =  12'b110101101000;     //371pi/512
   sin[372]  =  12'b110011111001;     //372pi/512
   cos[372]  =  12'b110101100011;     //372pi/512
   sin[373]  =  12'b110011111101;     //373pi/512
   cos[373]  =  12'b110101011110;     //373pi/512
   sin[374]  =  12'b110100000001;     //374pi/512
   cos[374]  =  12'b110101011010;     //374pi/512
   sin[375]  =  12'b110100000101;     //375pi/512
   cos[375]  =  12'b110101010101;     //375pi/512
   sin[376]  =  12'b110100001001;     //376pi/512
   cos[376]  =  12'b110101010000;     //376pi/512
   sin[377]  =  12'b110100001101;     //377pi/512
   cos[377]  =  12'b110101001100;     //377pi/512
   sin[378]  =  12'b110100010010;     //378pi/512
   cos[378]  =  12'b110101000111;     //378pi/512
   sin[379]  =  12'b110100010110;     //379pi/512
   cos[379]  =  12'b110101000010;     //379pi/512
   sin[380]  =  12'b110100011010;     //380pi/512
   cos[380]  =  12'b110100111110;     //380pi/512
   sin[381]  =  12'b110100011111;     //381pi/512
   cos[381]  =  12'b110100111001;     //381pi/512
   sin[382]  =  12'b110100100011;     //382pi/512
   cos[382]  =  12'b110100110101;     //382pi/512
   sin[383]  =  12'b110100100111;     //383pi/512
   cos[383]  =  12'b110100110000;     //383pi/512
   sin[384]  =  12'b110100101100;     //384pi/512
   cos[384]  =  12'b110100101100;     //384pi/512
   sin[385]  =  12'b110100110000;     //385pi/512
   cos[385]  =  12'b110100100111;     //385pi/512
   sin[386]  =  12'b110100110101;     //386pi/512
   cos[386]  =  12'b110100100011;     //386pi/512
   sin[387]  =  12'b110100111001;     //387pi/512
   cos[387]  =  12'b110100011111;     //387pi/512
   sin[388]  =  12'b110100111110;     //388pi/512
   cos[388]  =  12'b110100011010;     //388pi/512
   sin[389]  =  12'b110101000010;     //389pi/512
   cos[389]  =  12'b110100010110;     //389pi/512
   sin[390]  =  12'b110101000111;     //390pi/512
   cos[390]  =  12'b110100010010;     //390pi/512
   sin[391]  =  12'b110101001100;     //391pi/512
   cos[391]  =  12'b110100001101;     //391pi/512
   sin[392]  =  12'b110101010000;     //392pi/512
   cos[392]  =  12'b110100001001;     //392pi/512
   sin[393]  =  12'b110101010101;     //393pi/512
   cos[393]  =  12'b110100000101;     //393pi/512
   sin[394]  =  12'b110101011010;     //394pi/512
   cos[394]  =  12'b110100000001;     //394pi/512
   sin[395]  =  12'b110101011110;     //395pi/512
   cos[395]  =  12'b110011111101;     //395pi/512
   sin[396]  =  12'b110101100011;     //396pi/512
   cos[396]  =  12'b110011111001;     //396pi/512
   sin[397]  =  12'b110101101000;     //397pi/512
   cos[397]  =  12'b110011110101;     //397pi/512
   sin[398]  =  12'b110101101101;     //398pi/512
   cos[398]  =  12'b110011110000;     //398pi/512
   sin[399]  =  12'b110101110010;     //399pi/512
   cos[399]  =  12'b110011101100;     //399pi/512
   sin[400]  =  12'b110101110110;     //400pi/512
   cos[400]  =  12'b110011101000;     //400pi/512
   sin[401]  =  12'b110101111011;     //401pi/512
   cos[401]  =  12'b110011100100;     //401pi/512
   sin[402]  =  12'b110110000000;     //402pi/512
   cos[402]  =  12'b110011100001;     //402pi/512
   sin[403]  =  12'b110110000101;     //403pi/512
   cos[403]  =  12'b110011011101;     //403pi/512
   sin[404]  =  12'b110110001010;     //404pi/512
   cos[404]  =  12'b110011011001;     //404pi/512
   sin[405]  =  12'b110110001111;     //405pi/512
   cos[405]  =  12'b110011010101;     //405pi/512
   sin[406]  =  12'b110110010100;     //406pi/512
   cos[406]  =  12'b110011010001;     //406pi/512
   sin[407]  =  12'b110110011001;     //407pi/512
   cos[407]  =  12'b110011001101;     //407pi/512
   sin[408]  =  12'b110110011110;     //408pi/512
   cos[408]  =  12'b110011001010;     //408pi/512
   sin[409]  =  12'b110110100011;     //409pi/512
   cos[409]  =  12'b110011000110;     //409pi/512
   sin[410]  =  12'b110110101000;     //410pi/512
   cos[410]  =  12'b110011000010;     //410pi/512
   sin[411]  =  12'b110110101101;     //411pi/512
   cos[411]  =  12'b110010111110;     //411pi/512
   sin[412]  =  12'b110110110010;     //412pi/512
   cos[412]  =  12'b110010111011;     //412pi/512
   sin[413]  =  12'b110110111000;     //413pi/512
   cos[413]  =  12'b110010110111;     //413pi/512
   sin[414]  =  12'b110110111101;     //414pi/512
   cos[414]  =  12'b110010110100;     //414pi/512
   sin[415]  =  12'b110111000010;     //415pi/512
   cos[415]  =  12'b110010110000;     //415pi/512
   sin[416]  =  12'b110111000111;     //416pi/512
   cos[416]  =  12'b110010101101;     //416pi/512
   sin[417]  =  12'b110111001100;     //417pi/512
   cos[417]  =  12'b110010101001;     //417pi/512
   sin[418]  =  12'b110111010010;     //418pi/512
   cos[418]  =  12'b110010100110;     //418pi/512
   sin[419]  =  12'b110111010111;     //419pi/512
   cos[419]  =  12'b110010100010;     //419pi/512
   sin[420]  =  12'b110111011100;     //420pi/512
   cos[420]  =  12'b110010011111;     //420pi/512
   sin[421]  =  12'b110111100001;     //421pi/512
   cos[421]  =  12'b110010011100;     //421pi/512
   sin[422]  =  12'b110111100111;     //422pi/512
   cos[422]  =  12'b110010011000;     //422pi/512
   sin[423]  =  12'b110111101100;     //423pi/512
   cos[423]  =  12'b110010010101;     //423pi/512
   sin[424]  =  12'b110111110010;     //424pi/512
   cos[424]  =  12'b110010010010;     //424pi/512
   sin[425]  =  12'b110111110111;     //425pi/512
   cos[425]  =  12'b110010001110;     //425pi/512
   sin[426]  =  12'b110111111100;     //426pi/512
   cos[426]  =  12'b110010001011;     //426pi/512
   sin[427]  =  12'b111000000010;     //427pi/512
   cos[427]  =  12'b110010001000;     //427pi/512
   sin[428]  =  12'b111000000111;     //428pi/512
   cos[428]  =  12'b110010000101;     //428pi/512
   sin[429]  =  12'b111000001101;     //429pi/512
   cos[429]  =  12'b110010000010;     //429pi/512
   sin[430]  =  12'b111000010010;     //430pi/512
   cos[430]  =  12'b110001111111;     //430pi/512
   sin[431]  =  12'b111000011000;     //431pi/512
   cos[431]  =  12'b110001111100;     //431pi/512
   sin[432]  =  12'b111000011101;     //432pi/512
   cos[432]  =  12'b110001111001;     //432pi/512
   sin[433]  =  12'b111000100011;     //433pi/512
   cos[433]  =  12'b110001110110;     //433pi/512
   sin[434]  =  12'b111000101000;     //434pi/512
   cos[434]  =  12'b110001110011;     //434pi/512
   sin[435]  =  12'b111000101110;     //435pi/512
   cos[435]  =  12'b110001110000;     //435pi/512
   sin[436]  =  12'b111000110100;     //436pi/512
   cos[436]  =  12'b110001101101;     //436pi/512
   sin[437]  =  12'b111000111001;     //437pi/512
   cos[437]  =  12'b110001101011;     //437pi/512
   sin[438]  =  12'b111000111111;     //438pi/512
   cos[438]  =  12'b110001101000;     //438pi/512
   sin[439]  =  12'b111001000101;     //439pi/512
   cos[439]  =  12'b110001100101;     //439pi/512
   sin[440]  =  12'b111001001010;     //440pi/512
   cos[440]  =  12'b110001100010;     //440pi/512
   sin[441]  =  12'b111001010000;     //441pi/512
   cos[441]  =  12'b110001100000;     //441pi/512
   sin[442]  =  12'b111001010110;     //442pi/512
   cos[442]  =  12'b110001011101;     //442pi/512
   sin[443]  =  12'b111001011011;     //443pi/512
   cos[443]  =  12'b110001011010;     //443pi/512
   sin[444]  =  12'b111001100001;     //444pi/512
   cos[444]  =  12'b110001011000;     //444pi/512
   sin[445]  =  12'b111001100111;     //445pi/512
   cos[445]  =  12'b110001010101;     //445pi/512
   sin[446]  =  12'b111001101101;     //446pi/512
   cos[446]  =  12'b110001010011;     //446pi/512
   sin[447]  =  12'b111001110010;     //447pi/512
   cos[447]  =  12'b110001010000;     //447pi/512
   sin[448]  =  12'b111001111000;     //448pi/512
   cos[448]  =  12'b110001001110;     //448pi/512
   sin[449]  =  12'b111001111110;     //449pi/512
   cos[449]  =  12'b110001001100;     //449pi/512
   sin[450]  =  12'b111010000100;     //450pi/512
   cos[450]  =  12'b110001001001;     //450pi/512
   sin[451]  =  12'b111010001010;     //451pi/512
   cos[451]  =  12'b110001000111;     //451pi/512
   sin[452]  =  12'b111010001111;     //452pi/512
   cos[452]  =  12'b110001000101;     //452pi/512
   sin[453]  =  12'b111010010101;     //453pi/512
   cos[453]  =  12'b110001000010;     //453pi/512
   sin[454]  =  12'b111010011011;     //454pi/512
   cos[454]  =  12'b110001000000;     //454pi/512
   sin[455]  =  12'b111010100001;     //455pi/512
   cos[455]  =  12'b110000111110;     //455pi/512
   sin[456]  =  12'b111010100111;     //456pi/512
   cos[456]  =  12'b110000111100;     //456pi/512
   sin[457]  =  12'b111010101101;     //457pi/512
   cos[457]  =  12'b110000111010;     //457pi/512
   sin[458]  =  12'b111010110011;     //458pi/512
   cos[458]  =  12'b110000111000;     //458pi/512
   sin[459]  =  12'b111010111001;     //459pi/512
   cos[459]  =  12'b110000110110;     //459pi/512
   sin[460]  =  12'b111010111111;     //460pi/512
   cos[460]  =  12'b110000110100;     //460pi/512
   sin[461]  =  12'b111011000101;     //461pi/512
   cos[461]  =  12'b110000110010;     //461pi/512
   sin[462]  =  12'b111011001011;     //462pi/512
   cos[462]  =  12'b110000110000;     //462pi/512
   sin[463]  =  12'b111011010001;     //463pi/512
   cos[463]  =  12'b110000101110;     //463pi/512
   sin[464]  =  12'b111011010111;     //464pi/512
   cos[464]  =  12'b110000101100;     //464pi/512
   sin[465]  =  12'b111011011101;     //465pi/512
   cos[465]  =  12'b110000101010;     //465pi/512
   sin[466]  =  12'b111011100011;     //466pi/512
   cos[466]  =  12'b110000101001;     //466pi/512
   sin[467]  =  12'b111011101001;     //467pi/512
   cos[467]  =  12'b110000100111;     //467pi/512
   sin[468]  =  12'b111011101111;     //468pi/512
   cos[468]  =  12'b110000100101;     //468pi/512
   sin[469]  =  12'b111011110101;     //469pi/512
   cos[469]  =  12'b110000100011;     //469pi/512
   sin[470]  =  12'b111011111011;     //470pi/512
   cos[470]  =  12'b110000100010;     //470pi/512
   sin[471]  =  12'b111100000001;     //471pi/512
   cos[471]  =  12'b110000100000;     //471pi/512
   sin[472]  =  12'b111100000111;     //472pi/512
   cos[472]  =  12'b110000011111;     //472pi/512
   sin[473]  =  12'b111100001101;     //473pi/512
   cos[473]  =  12'b110000011101;     //473pi/512
   sin[474]  =  12'b111100010011;     //474pi/512
   cos[474]  =  12'b110000011100;     //474pi/512
   sin[475]  =  12'b111100011010;     //475pi/512
   cos[475]  =  12'b110000011010;     //475pi/512
   sin[476]  =  12'b111100100000;     //476pi/512
   cos[476]  =  12'b110000011001;     //476pi/512
   sin[477]  =  12'b111100100110;     //477pi/512
   cos[477]  =  12'b110000011000;     //477pi/512
   sin[478]  =  12'b111100101100;     //478pi/512
   cos[478]  =  12'b110000010110;     //478pi/512
   sin[479]  =  12'b111100110010;     //479pi/512
   cos[479]  =  12'b110000010101;     //479pi/512
   sin[480]  =  12'b111100111000;     //480pi/512
   cos[480]  =  12'b110000010100;     //480pi/512
   sin[481]  =  12'b111100111110;     //481pi/512
   cos[481]  =  12'b110000010010;     //481pi/512
   sin[482]  =  12'b111101000101;     //482pi/512
   cos[482]  =  12'b110000010001;     //482pi/512
   sin[483]  =  12'b111101001011;     //483pi/512
   cos[483]  =  12'b110000010000;     //483pi/512
   sin[484]  =  12'b111101010001;     //484pi/512
   cos[484]  =  12'b110000001111;     //484pi/512
   sin[485]  =  12'b111101010111;     //485pi/512
   cos[485]  =  12'b110000001110;     //485pi/512
   sin[486]  =  12'b111101011101;     //486pi/512
   cos[486]  =  12'b110000001101;     //486pi/512
   sin[487]  =  12'b111101100100;     //487pi/512
   cos[487]  =  12'b110000001100;     //487pi/512
   sin[488]  =  12'b111101101010;     //488pi/512
   cos[488]  =  12'b110000001011;     //488pi/512
   sin[489]  =  12'b111101110000;     //489pi/512
   cos[489]  =  12'b110000001010;     //489pi/512
   sin[490]  =  12'b111101110110;     //490pi/512
   cos[490]  =  12'b110000001001;     //490pi/512
   sin[491]  =  12'b111101111100;     //491pi/512
   cos[491]  =  12'b110000001000;     //491pi/512
   sin[492]  =  12'b111110000011;     //492pi/512
   cos[492]  =  12'b110000001000;     //492pi/512
   sin[493]  =  12'b111110001001;     //493pi/512
   cos[493]  =  12'b110000000111;     //493pi/512
   sin[494]  =  12'b111110001111;     //494pi/512
   cos[494]  =  12'b110000000110;     //494pi/512
   sin[495]  =  12'b111110010101;     //495pi/512
   cos[495]  =  12'b110000000110;     //495pi/512
   sin[496]  =  12'b111110011100;     //496pi/512
   cos[496]  =  12'b110000000101;     //496pi/512
   sin[497]  =  12'b111110100010;     //497pi/512
   cos[497]  =  12'b110000000100;     //497pi/512
   sin[498]  =  12'b111110101000;     //498pi/512
   cos[498]  =  12'b110000000100;     //498pi/512
   sin[499]  =  12'b111110101110;     //499pi/512
   cos[499]  =  12'b110000000011;     //499pi/512
   sin[500]  =  12'b111110110101;     //500pi/512
   cos[500]  =  12'b110000000011;     //500pi/512
   sin[501]  =  12'b111110111011;     //501pi/512
   cos[501]  =  12'b110000000010;     //501pi/512
   sin[502]  =  12'b111111000001;     //502pi/512
   cos[502]  =  12'b110000000010;     //502pi/512
   sin[503]  =  12'b111111000111;     //503pi/512
   cos[503]  =  12'b110000000010;     //503pi/512
   sin[504]  =  12'b111111001110;     //504pi/512
   cos[504]  =  12'b110000000001;     //504pi/512
   sin[505]  =  12'b111111010100;     //505pi/512
   cos[505]  =  12'b110000000001;     //505pi/512
   sin[506]  =  12'b111111011010;     //506pi/512
   cos[506]  =  12'b110000000001;     //506pi/512
   sin[507]  =  12'b111111100001;     //507pi/512
   cos[507]  =  12'b110000000000;     //507pi/512
   sin[508]  =  12'b111111100111;     //508pi/512
   cos[508]  =  12'b110000000000;     //508pi/512
   sin[509]  =  12'b111111101101;     //509pi/512
   cos[509]  =  12'b110000000000;     //509pi/512
   sin[510]  =  12'b111111110011;     //510pi/512
   cos[510]  =  12'b110000000000;     //510pi/512
   sin[511]  =  12'b111111111010;     //511pi/512
   cos[511]  =  12'b110000000000;     //511pi/512
   m_sin[0]  =  12'b000000000000;     //0pi/512
   m_cos[0]  =  12'b010000000000;     //0pi/512
   m_sin[1]  =  12'b111111111010;     //1pi/512
   m_cos[1]  =  12'b001111111111;     //1pi/512
   m_sin[2]  =  12'b111111110101;     //2pi/512
   m_cos[2]  =  12'b001111111111;     //2pi/512
   m_sin[3]  =  12'b111111101111;     //3pi/512
   m_cos[3]  =  12'b001111111111;     //3pi/512
   m_sin[4]  =  12'b111111101001;     //4pi/512
   m_cos[4]  =  12'b001111111111;     //4pi/512
   m_sin[5]  =  12'b111111100100;     //5pi/512
   m_cos[5]  =  12'b001111111111;     //5pi/512
   m_sin[6]  =  12'b111111011110;     //6pi/512
   m_cos[6]  =  12'b001111111111;     //6pi/512
   m_sin[7]  =  12'b111111011000;     //7pi/512
   m_cos[7]  =  12'b001111111111;     //7pi/512
   m_sin[8]  =  12'b111111010011;     //8pi/512
   m_cos[8]  =  12'b001111111111;     //8pi/512
   m_sin[9]  =  12'b111111001101;     //9pi/512
   m_cos[9]  =  12'b001111111110;     //9pi/512
   m_sin[10]  =  12'b111111000111;     //10pi/512
   m_cos[10]  =  12'b001111111110;     //10pi/512
   m_sin[11]  =  12'b111111000010;     //11pi/512
   m_cos[11]  =  12'b001111111110;     //11pi/512
   m_sin[12]  =  12'b111110111100;     //12pi/512
   m_cos[12]  =  12'b001111111101;     //12pi/512
   m_sin[13]  =  12'b111110110111;     //13pi/512
   m_cos[13]  =  12'b001111111101;     //13pi/512
   m_sin[14]  =  12'b111110110001;     //14pi/512
   m_cos[14]  =  12'b001111111100;     //14pi/512
   m_sin[15]  =  12'b111110101011;     //15pi/512
   m_cos[15]  =  12'b001111111100;     //15pi/512
   m_sin[16]  =  12'b111110100110;     //16pi/512
   m_cos[16]  =  12'b001111111100;     //16pi/512
   m_sin[17]  =  12'b111110100000;     //17pi/512
   m_cos[17]  =  12'b001111111011;     //17pi/512
   m_sin[18]  =  12'b111110011010;     //18pi/512
   m_cos[18]  =  12'b001111111010;     //18pi/512
   m_sin[19]  =  12'b111110010101;     //19pi/512
   m_cos[19]  =  12'b001111111010;     //19pi/512
   m_sin[20]  =  12'b111110001111;     //20pi/512
   m_cos[20]  =  12'b001111111001;     //20pi/512
   m_sin[21]  =  12'b111110001010;     //21pi/512
   m_cos[21]  =  12'b001111111001;     //21pi/512
   m_sin[22]  =  12'b111110000100;     //22pi/512
   m_cos[22]  =  12'b001111111000;     //22pi/512
   m_sin[23]  =  12'b111101111110;     //23pi/512
   m_cos[23]  =  12'b001111110111;     //23pi/512
   m_sin[24]  =  12'b111101111001;     //24pi/512
   m_cos[24]  =  12'b001111110111;     //24pi/512
   m_sin[25]  =  12'b111101110011;     //25pi/512
   m_cos[25]  =  12'b001111110110;     //25pi/512
   m_sin[26]  =  12'b111101101101;     //26pi/512
   m_cos[26]  =  12'b001111110101;     //26pi/512
   m_sin[27]  =  12'b111101101000;     //27pi/512
   m_cos[27]  =  12'b001111110100;     //27pi/512
   m_sin[28]  =  12'b111101100010;     //28pi/512
   m_cos[28]  =  12'b001111110011;     //28pi/512
   m_sin[29]  =  12'b111101011101;     //29pi/512
   m_cos[29]  =  12'b001111110010;     //29pi/512
   m_sin[30]  =  12'b111101010111;     //30pi/512
   m_cos[30]  =  12'b001111110001;     //30pi/512
   m_sin[31]  =  12'b111101010010;     //31pi/512
   m_cos[31]  =  12'b001111110001;     //31pi/512
   m_sin[32]  =  12'b111101001100;     //32pi/512
   m_cos[32]  =  12'b001111110000;     //32pi/512
   m_sin[33]  =  12'b111101000110;     //33pi/512
   m_cos[33]  =  12'b001111101111;     //33pi/512
   m_sin[34]  =  12'b111101000001;     //34pi/512
   m_cos[34]  =  12'b001111101110;     //34pi/512
   m_sin[35]  =  12'b111100111011;     //35pi/512
   m_cos[35]  =  12'b001111101100;     //35pi/512
   m_sin[36]  =  12'b111100110110;     //36pi/512
   m_cos[36]  =  12'b001111101011;     //36pi/512
   m_sin[37]  =  12'b111100110000;     //37pi/512
   m_cos[37]  =  12'b001111101010;     //37pi/512
   m_sin[38]  =  12'b111100101011;     //38pi/512
   m_cos[38]  =  12'b001111101001;     //38pi/512
   m_sin[39]  =  12'b111100100101;     //39pi/512
   m_cos[39]  =  12'b001111101000;     //39pi/512
   m_sin[40]  =  12'b111100100000;     //40pi/512
   m_cos[40]  =  12'b001111100111;     //40pi/512
   m_sin[41]  =  12'b111100011010;     //41pi/512
   m_cos[41]  =  12'b001111100101;     //41pi/512
   m_sin[42]  =  12'b111100010101;     //42pi/512
   m_cos[42]  =  12'b001111100100;     //42pi/512
   m_sin[43]  =  12'b111100001111;     //43pi/512
   m_cos[43]  =  12'b001111100011;     //43pi/512
   m_sin[44]  =  12'b111100001010;     //44pi/512
   m_cos[44]  =  12'b001111100001;     //44pi/512
   m_sin[45]  =  12'b111100000100;     //45pi/512
   m_cos[45]  =  12'b001111100000;     //45pi/512
   m_sin[46]  =  12'b111011111111;     //46pi/512
   m_cos[46]  =  12'b001111011111;     //46pi/512
   m_sin[47]  =  12'b111011111001;     //47pi/512
   m_cos[47]  =  12'b001111011101;     //47pi/512
   m_sin[48]  =  12'b111011110100;     //48pi/512
   m_cos[48]  =  12'b001111011100;     //48pi/512
   m_sin[49]  =  12'b111011101110;     //49pi/512
   m_cos[49]  =  12'b001111011010;     //49pi/512
   m_sin[50]  =  12'b111011101001;     //50pi/512
   m_cos[50]  =  12'b001111011001;     //50pi/512
   m_sin[51]  =  12'b111011100011;     //51pi/512
   m_cos[51]  =  12'b001111010111;     //51pi/512
   m_sin[52]  =  12'b111011011110;     //52pi/512
   m_cos[52]  =  12'b001111010110;     //52pi/512
   m_sin[53]  =  12'b111011011001;     //53pi/512
   m_cos[53]  =  12'b001111010100;     //53pi/512
   m_sin[54]  =  12'b111011010011;     //54pi/512
   m_cos[54]  =  12'b001111010010;     //54pi/512
   m_sin[55]  =  12'b111011001110;     //55pi/512
   m_cos[55]  =  12'b001111010001;     //55pi/512
   m_sin[56]  =  12'b111011001000;     //56pi/512
   m_cos[56]  =  12'b001111001111;     //56pi/512
   m_sin[57]  =  12'b111011000011;     //57pi/512
   m_cos[57]  =  12'b001111001101;     //57pi/512
   m_sin[58]  =  12'b111010111110;     //58pi/512
   m_cos[58]  =  12'b001111001011;     //58pi/512
   m_sin[59]  =  12'b111010111000;     //59pi/512
   m_cos[59]  =  12'b001111001010;     //59pi/512
   m_sin[60]  =  12'b111010110011;     //60pi/512
   m_cos[60]  =  12'b001111001000;     //60pi/512
   m_sin[61]  =  12'b111010101110;     //61pi/512
   m_cos[61]  =  12'b001111000110;     //61pi/512
   m_sin[62]  =  12'b111010101000;     //62pi/512
   m_cos[62]  =  12'b001111000100;     //62pi/512
   m_sin[63]  =  12'b111010100011;     //63pi/512
   m_cos[63]  =  12'b001111000010;     //63pi/512
   m_sin[64]  =  12'b111010011110;     //64pi/512
   m_cos[64]  =  12'b001111000000;     //64pi/512
   m_sin[65]  =  12'b111010011000;     //65pi/512
   m_cos[65]  =  12'b001110111110;     //65pi/512
   m_sin[66]  =  12'b111010010011;     //66pi/512
   m_cos[66]  =  12'b001110111100;     //66pi/512
   m_sin[67]  =  12'b111010001110;     //67pi/512
   m_cos[67]  =  12'b001110111010;     //67pi/512
   m_sin[68]  =  12'b111010001000;     //68pi/512
   m_cos[68]  =  12'b001110111000;     //68pi/512
   m_sin[69]  =  12'b111010000011;     //69pi/512
   m_cos[69]  =  12'b001110110110;     //69pi/512
   m_sin[70]  =  12'b111001111110;     //70pi/512
   m_cos[70]  =  12'b001110110100;     //70pi/512
   m_sin[71]  =  12'b111001111001;     //71pi/512
   m_cos[71]  =  12'b001110110010;     //71pi/512
   m_sin[72]  =  12'b111001110011;     //72pi/512
   m_cos[72]  =  12'b001110110000;     //72pi/512
   m_sin[73]  =  12'b111001101110;     //73pi/512
   m_cos[73]  =  12'b001110101101;     //73pi/512
   m_sin[74]  =  12'b111001101001;     //74pi/512
   m_cos[74]  =  12'b001110101011;     //74pi/512
   m_sin[75]  =  12'b111001100100;     //75pi/512
   m_cos[75]  =  12'b001110101001;     //75pi/512
   m_sin[76]  =  12'b111001011111;     //76pi/512
   m_cos[76]  =  12'b001110100111;     //76pi/512
   m_sin[77]  =  12'b111001011010;     //77pi/512
   m_cos[77]  =  12'b001110100100;     //77pi/512
   m_sin[78]  =  12'b111001010100;     //78pi/512
   m_cos[78]  =  12'b001110100010;     //78pi/512
   m_sin[79]  =  12'b111001001111;     //79pi/512
   m_cos[79]  =  12'b001110100000;     //79pi/512
   m_sin[80]  =  12'b111001001010;     //80pi/512
   m_cos[80]  =  12'b001110011101;     //80pi/512
   m_sin[81]  =  12'b111001000101;     //81pi/512
   m_cos[81]  =  12'b001110011011;     //81pi/512
   m_sin[82]  =  12'b111001000000;     //82pi/512
   m_cos[82]  =  12'b001110011000;     //82pi/512
   m_sin[83]  =  12'b111000111011;     //83pi/512
   m_cos[83]  =  12'b001110010110;     //83pi/512
   m_sin[84]  =  12'b111000110110;     //84pi/512
   m_cos[84]  =  12'b001110010011;     //84pi/512
   m_sin[85]  =  12'b111000110001;     //85pi/512
   m_cos[85]  =  12'b001110010001;     //85pi/512
   m_sin[86]  =  12'b111000101100;     //86pi/512
   m_cos[86]  =  12'b001110001110;     //86pi/512
   m_sin[87]  =  12'b111000100111;     //87pi/512
   m_cos[87]  =  12'b001110001100;     //87pi/512
   m_sin[88]  =  12'b111000100010;     //88pi/512
   m_cos[88]  =  12'b001110001001;     //88pi/512
   m_sin[89]  =  12'b111000011101;     //89pi/512
   m_cos[89]  =  12'b001110000110;     //89pi/512
   m_sin[90]  =  12'b111000011000;     //90pi/512
   m_cos[90]  =  12'b001110000100;     //90pi/512
   m_sin[91]  =  12'b111000010011;     //91pi/512
   m_cos[91]  =  12'b001110000001;     //91pi/512
   m_sin[92]  =  12'b111000001110;     //92pi/512
   m_cos[92]  =  12'b001101111110;     //92pi/512
   m_sin[93]  =  12'b111000001001;     //93pi/512
   m_cos[93]  =  12'b001101111011;     //93pi/512
   m_sin[94]  =  12'b111000000100;     //94pi/512
   m_cos[94]  =  12'b001101111001;     //94pi/512
   m_sin[95]  =  12'b110111111111;     //95pi/512
   m_cos[95]  =  12'b001101110110;     //95pi/512
   m_sin[96]  =  12'b110111111010;     //96pi/512
   m_cos[96]  =  12'b001101110011;     //96pi/512
   m_sin[97]  =  12'b110111110101;     //97pi/512
   m_cos[97]  =  12'b001101110000;     //97pi/512
   m_sin[98]  =  12'b110111110000;     //98pi/512
   m_cos[98]  =  12'b001101101101;     //98pi/512
   m_sin[99]  =  12'b110111101100;     //99pi/512
   m_cos[99]  =  12'b001101101010;     //99pi/512
   m_sin[100]  =  12'b110111100111;     //100pi/512
   m_cos[100]  =  12'b001101100111;     //100pi/512
   m_sin[101]  =  12'b110111100010;     //101pi/512
   m_cos[101]  =  12'b001101100100;     //101pi/512
   m_sin[102]  =  12'b110111011101;     //102pi/512
   m_cos[102]  =  12'b001101100001;     //102pi/512
   m_sin[103]  =  12'b110111011000;     //103pi/512
   m_cos[103]  =  12'b001101011110;     //103pi/512
   m_sin[104]  =  12'b110111010100;     //104pi/512
   m_cos[104]  =  12'b001101011011;     //104pi/512
   m_sin[105]  =  12'b110111001111;     //105pi/512
   m_cos[105]  =  12'b001101011000;     //105pi/512
   m_sin[106]  =  12'b110111001010;     //106pi/512
   m_cos[106]  =  12'b001101010101;     //106pi/512
   m_sin[107]  =  12'b110111000110;     //107pi/512
   m_cos[107]  =  12'b001101010010;     //107pi/512
   m_sin[108]  =  12'b110111000001;     //108pi/512
   m_cos[108]  =  12'b001101001111;     //108pi/512
   m_sin[109]  =  12'b110110111100;     //109pi/512
   m_cos[109]  =  12'b001101001100;     //109pi/512
   m_sin[110]  =  12'b110110111000;     //110pi/512
   m_cos[110]  =  12'b001101001000;     //110pi/512
   m_sin[111]  =  12'b110110110011;     //111pi/512
   m_cos[111]  =  12'b001101000101;     //111pi/512
   m_sin[112]  =  12'b110110101110;     //112pi/512
   m_cos[112]  =  12'b001101000010;     //112pi/512
   m_sin[113]  =  12'b110110101010;     //113pi/512
   m_cos[113]  =  12'b001100111111;     //113pi/512
   m_sin[114]  =  12'b110110100101;     //114pi/512
   m_cos[114]  =  12'b001100111011;     //114pi/512
   m_sin[115]  =  12'b110110100001;     //115pi/512
   m_cos[115]  =  12'b001100111000;     //115pi/512
   m_sin[116]  =  12'b110110011100;     //116pi/512
   m_cos[116]  =  12'b001100110100;     //116pi/512
   m_sin[117]  =  12'b110110010111;     //117pi/512
   m_cos[117]  =  12'b001100110001;     //117pi/512
   m_sin[118]  =  12'b110110010011;     //118pi/512
   m_cos[118]  =  12'b001100101110;     //118pi/512
   m_sin[119]  =  12'b110110001110;     //119pi/512
   m_cos[119]  =  12'b001100101010;     //119pi/512
   m_sin[120]  =  12'b110110001010;     //120pi/512
   m_cos[120]  =  12'b001100100111;     //120pi/512
   m_sin[121]  =  12'b110110000110;     //121pi/512
   m_cos[121]  =  12'b001100100011;     //121pi/512
   m_sin[122]  =  12'b110110000001;     //122pi/512
   m_cos[122]  =  12'b001100100000;     //122pi/512
   m_sin[123]  =  12'b110101111101;     //123pi/512
   m_cos[123]  =  12'b001100011100;     //123pi/512
   m_sin[124]  =  12'b110101111000;     //124pi/512
   m_cos[124]  =  12'b001100011001;     //124pi/512
   m_sin[125]  =  12'b110101110100;     //125pi/512
   m_cos[125]  =  12'b001100010101;     //125pi/512
   m_sin[126]  =  12'b110101110000;     //126pi/512
   m_cos[126]  =  12'b001100010001;     //126pi/512
   m_sin[127]  =  12'b110101101011;     //127pi/512
   m_cos[127]  =  12'b001100001110;     //127pi/512
   m_sin[128]  =  12'b110101100111;     //128pi/512
   m_cos[128]  =  12'b001100001010;     //128pi/512
   m_sin[129]  =  12'b110101100011;     //129pi/512
   m_cos[129]  =  12'b001100000110;     //129pi/512
   m_sin[130]  =  12'b110101011110;     //130pi/512
   m_cos[130]  =  12'b001100000011;     //130pi/512
   m_sin[131]  =  12'b110101011010;     //131pi/512
   m_cos[131]  =  12'b001011111111;     //131pi/512
   m_sin[132]  =  12'b110101010110;     //132pi/512
   m_cos[132]  =  12'b001011111011;     //132pi/512
   m_sin[133]  =  12'b110101010010;     //133pi/512
   m_cos[133]  =  12'b001011110111;     //133pi/512
   m_sin[134]  =  12'b110101001110;     //134pi/512
   m_cos[134]  =  12'b001011110100;     //134pi/512
   m_sin[135]  =  12'b110101001001;     //135pi/512
   m_cos[135]  =  12'b001011110000;     //135pi/512
   m_sin[136]  =  12'b110101000101;     //136pi/512
   m_cos[136]  =  12'b001011101100;     //136pi/512
   m_sin[137]  =  12'b110101000001;     //137pi/512
   m_cos[137]  =  12'b001011101000;     //137pi/512
   m_sin[138]  =  12'b110100111101;     //138pi/512
   m_cos[138]  =  12'b001011100100;     //138pi/512
   m_sin[139]  =  12'b110100111001;     //139pi/512
   m_cos[139]  =  12'b001011100000;     //139pi/512
   m_sin[140]  =  12'b110100110101;     //140pi/512
   m_cos[140]  =  12'b001011011100;     //140pi/512
   m_sin[141]  =  12'b110100110001;     //141pi/512
   m_cos[141]  =  12'b001011011000;     //141pi/512
   m_sin[142]  =  12'b110100101101;     //142pi/512
   m_cos[142]  =  12'b001011010100;     //142pi/512
   m_sin[143]  =  12'b110100101001;     //143pi/512
   m_cos[143]  =  12'b001011010000;     //143pi/512
   m_sin[144]  =  12'b110100100101;     //144pi/512
   m_cos[144]  =  12'b001011001100;     //144pi/512
   m_sin[145]  =  12'b110100100001;     //145pi/512
   m_cos[145]  =  12'b001011001000;     //145pi/512
   m_sin[146]  =  12'b110100011101;     //146pi/512
   m_cos[146]  =  12'b001011000100;     //146pi/512
   m_sin[147]  =  12'b110100011001;     //147pi/512
   m_cos[147]  =  12'b001011000000;     //147pi/512
   m_sin[148]  =  12'b110100010101;     //148pi/512
   m_cos[148]  =  12'b001010111100;     //148pi/512
   m_sin[149]  =  12'b110100010001;     //149pi/512
   m_cos[149]  =  12'b001010111000;     //149pi/512
   m_sin[150]  =  12'b110100001101;     //150pi/512
   m_cos[150]  =  12'b001010110100;     //150pi/512
   m_sin[151]  =  12'b110100001010;     //151pi/512
   m_cos[151]  =  12'b001010110000;     //151pi/512
   m_sin[152]  =  12'b110100000110;     //152pi/512
   m_cos[152]  =  12'b001010101011;     //152pi/512
   m_sin[153]  =  12'b110100000010;     //153pi/512
   m_cos[153]  =  12'b001010100111;     //153pi/512
   m_sin[154]  =  12'b110011111110;     //154pi/512
   m_cos[154]  =  12'b001010100011;     //154pi/512
   m_sin[155]  =  12'b110011111011;     //155pi/512
   m_cos[155]  =  12'b001010011111;     //155pi/512
   m_sin[156]  =  12'b110011110111;     //156pi/512
   m_cos[156]  =  12'b001010011010;     //156pi/512
   m_sin[157]  =  12'b110011110011;     //157pi/512
   m_cos[157]  =  12'b001010010110;     //157pi/512
   m_sin[158]  =  12'b110011110000;     //158pi/512
   m_cos[158]  =  12'b001010010010;     //158pi/512
   m_sin[159]  =  12'b110011101100;     //159pi/512
   m_cos[159]  =  12'b001010001101;     //159pi/512
   m_sin[160]  =  12'b110011101000;     //160pi/512
   m_cos[160]  =  12'b001010001001;     //160pi/512
   m_sin[161]  =  12'b110011100101;     //161pi/512
   m_cos[161]  =  12'b001010000101;     //161pi/512
   m_sin[162]  =  12'b110011100001;     //162pi/512
   m_cos[162]  =  12'b001010000000;     //162pi/512
   m_sin[163]  =  12'b110011011110;     //163pi/512
   m_cos[163]  =  12'b001001111100;     //163pi/512
   m_sin[164]  =  12'b110011011010;     //164pi/512
   m_cos[164]  =  12'b001001110111;     //164pi/512
   m_sin[165]  =  12'b110011010111;     //165pi/512
   m_cos[165]  =  12'b001001110011;     //165pi/512
   m_sin[166]  =  12'b110011010011;     //166pi/512
   m_cos[166]  =  12'b001001101111;     //166pi/512
   m_sin[167]  =  12'b110011010000;     //167pi/512
   m_cos[167]  =  12'b001001101010;     //167pi/512
   m_sin[168]  =  12'b110011001101;     //168pi/512
   m_cos[168]  =  12'b001001100110;     //168pi/512
   m_sin[169]  =  12'b110011001001;     //169pi/512
   m_cos[169]  =  12'b001001100001;     //169pi/512
   m_sin[170]  =  12'b110011000110;     //170pi/512
   m_cos[170]  =  12'b001001011100;     //170pi/512
   m_sin[171]  =  12'b110011000010;     //171pi/512
   m_cos[171]  =  12'b001001011000;     //171pi/512
   m_sin[172]  =  12'b110010111111;     //172pi/512
   m_cos[172]  =  12'b001001010011;     //172pi/512
   m_sin[173]  =  12'b110010111100;     //173pi/512
   m_cos[173]  =  12'b001001001111;     //173pi/512
   m_sin[174]  =  12'b110010111001;     //174pi/512
   m_cos[174]  =  12'b001001001010;     //174pi/512
   m_sin[175]  =  12'b110010110101;     //175pi/512
   m_cos[175]  =  12'b001001000101;     //175pi/512
   m_sin[176]  =  12'b110010110010;     //176pi/512
   m_cos[176]  =  12'b001001000001;     //176pi/512
   m_sin[177]  =  12'b110010101111;     //177pi/512
   m_cos[177]  =  12'b001000111100;     //177pi/512
   m_sin[178]  =  12'b110010101100;     //178pi/512
   m_cos[178]  =  12'b001000110111;     //178pi/512
   m_sin[179]  =  12'b110010101001;     //179pi/512
   m_cos[179]  =  12'b001000110011;     //179pi/512
   m_sin[180]  =  12'b110010100110;     //180pi/512
   m_cos[180]  =  12'b001000101110;     //180pi/512
   m_sin[181]  =  12'b110010100011;     //181pi/512
   m_cos[181]  =  12'b001000101001;     //181pi/512
   m_sin[182]  =  12'b110010100000;     //182pi/512
   m_cos[182]  =  12'b001000100100;     //182pi/512
   m_sin[183]  =  12'b110010011101;     //183pi/512
   m_cos[183]  =  12'b001000100000;     //183pi/512
   m_sin[184]  =  12'b110010011010;     //184pi/512
   m_cos[184]  =  12'b001000011011;     //184pi/512
   m_sin[185]  =  12'b110010010111;     //185pi/512
   m_cos[185]  =  12'b001000010110;     //185pi/512
   m_sin[186]  =  12'b110010010100;     //186pi/512
   m_cos[186]  =  12'b001000010001;     //186pi/512
   m_sin[187]  =  12'b110010010001;     //187pi/512
   m_cos[187]  =  12'b001000001100;     //187pi/512
   m_sin[188]  =  12'b110010001110;     //188pi/512
   m_cos[188]  =  12'b001000000111;     //188pi/512
   m_sin[189]  =  12'b110010001011;     //189pi/512
   m_cos[189]  =  12'b001000000011;     //189pi/512
   m_sin[190]  =  12'b110010001000;     //190pi/512
   m_cos[190]  =  12'b000111111110;     //190pi/512
   m_sin[191]  =  12'b110010000101;     //191pi/512
   m_cos[191]  =  12'b000111111001;     //191pi/512
   m_sin[192]  =  12'b110010000011;     //192pi/512
   m_cos[192]  =  12'b000111110100;     //192pi/512
   m_sin[193]  =  12'b110010000000;     //193pi/512
   m_cos[193]  =  12'b000111101111;     //193pi/512
   m_sin[194]  =  12'b110001111101;     //194pi/512
   m_cos[194]  =  12'b000111101010;     //194pi/512
   m_sin[195]  =  12'b110001111010;     //195pi/512
   m_cos[195]  =  12'b000111100101;     //195pi/512
   m_sin[196]  =  12'b110001111000;     //196pi/512
   m_cos[196]  =  12'b000111100000;     //196pi/512
   m_sin[197]  =  12'b110001110101;     //197pi/512
   m_cos[197]  =  12'b000111011011;     //197pi/512
   m_sin[198]  =  12'b110001110010;     //198pi/512
   m_cos[198]  =  12'b000111010110;     //198pi/512
   m_sin[199]  =  12'b110001110000;     //199pi/512
   m_cos[199]  =  12'b000111010001;     //199pi/512
   m_sin[200]  =  12'b110001101101;     //200pi/512
   m_cos[200]  =  12'b000111001100;     //200pi/512
   m_sin[201]  =  12'b110001101011;     //201pi/512
   m_cos[201]  =  12'b000111000111;     //201pi/512
   m_sin[202]  =  12'b110001101000;     //202pi/512
   m_cos[202]  =  12'b000111000010;     //202pi/512
   m_sin[203]  =  12'b110001100110;     //203pi/512
   m_cos[203]  =  12'b000110111101;     //203pi/512
   m_sin[204]  =  12'b110001100011;     //204pi/512
   m_cos[204]  =  12'b000110111000;     //204pi/512
   m_sin[205]  =  12'b110001100001;     //205pi/512
   m_cos[205]  =  12'b000110110010;     //205pi/512
   m_sin[206]  =  12'b110001011111;     //206pi/512
   m_cos[206]  =  12'b000110101101;     //206pi/512
   m_sin[207]  =  12'b110001011100;     //207pi/512
   m_cos[207]  =  12'b000110101000;     //207pi/512
   m_sin[208]  =  12'b110001011010;     //208pi/512
   m_cos[208]  =  12'b000110100011;     //208pi/512
   m_sin[209]  =  12'b110001011000;     //209pi/512
   m_cos[209]  =  12'b000110011110;     //209pi/512
   m_sin[210]  =  12'b110001010101;     //210pi/512
   m_cos[210]  =  12'b000110011001;     //210pi/512
   m_sin[211]  =  12'b110001010011;     //211pi/512
   m_cos[211]  =  12'b000110010100;     //211pi/512
   m_sin[212]  =  12'b110001010001;     //212pi/512
   m_cos[212]  =  12'b000110001110;     //212pi/512
   m_sin[213]  =  12'b110001001111;     //213pi/512
   m_cos[213]  =  12'b000110001001;     //213pi/512
   m_sin[214]  =  12'b110001001101;     //214pi/512
   m_cos[214]  =  12'b000110000100;     //214pi/512
   m_sin[215]  =  12'b110001001010;     //215pi/512
   m_cos[215]  =  12'b000101111111;     //215pi/512
   m_sin[216]  =  12'b110001001000;     //216pi/512
   m_cos[216]  =  12'b000101111001;     //216pi/512
   m_sin[217]  =  12'b110001000110;     //217pi/512
   m_cos[217]  =  12'b000101110100;     //217pi/512
   m_sin[218]  =  12'b110001000100;     //218pi/512
   m_cos[218]  =  12'b000101101111;     //218pi/512
   m_sin[219]  =  12'b110001000010;     //219pi/512
   m_cos[219]  =  12'b000101101010;     //219pi/512
   m_sin[220]  =  12'b110001000000;     //220pi/512
   m_cos[220]  =  12'b000101100100;     //220pi/512
   m_sin[221]  =  12'b110000111110;     //221pi/512
   m_cos[221]  =  12'b000101011111;     //221pi/512
   m_sin[222]  =  12'b110000111100;     //222pi/512
   m_cos[222]  =  12'b000101011010;     //222pi/512
   m_sin[223]  =  12'b110000111010;     //223pi/512
   m_cos[223]  =  12'b000101010100;     //223pi/512
   m_sin[224]  =  12'b110000111001;     //224pi/512
   m_cos[224]  =  12'b000101001111;     //224pi/512
   m_sin[225]  =  12'b110000110111;     //225pi/512
   m_cos[225]  =  12'b000101001010;     //225pi/512
   m_sin[226]  =  12'b110000110101;     //226pi/512
   m_cos[226]  =  12'b000101000100;     //226pi/512
   m_sin[227]  =  12'b110000110011;     //227pi/512
   m_cos[227]  =  12'b000100111111;     //227pi/512
   m_sin[228]  =  12'b110000110001;     //228pi/512
   m_cos[228]  =  12'b000100111010;     //228pi/512
   m_sin[229]  =  12'b110000110000;     //229pi/512
   m_cos[229]  =  12'b000100110100;     //229pi/512
   m_sin[230]  =  12'b110000101110;     //230pi/512
   m_cos[230]  =  12'b000100101111;     //230pi/512
   m_sin[231]  =  12'b110000101100;     //231pi/512
   m_cos[231]  =  12'b000100101001;     //231pi/512
   m_sin[232]  =  12'b110000101011;     //232pi/512
   m_cos[232]  =  12'b000100100100;     //232pi/512
   m_sin[233]  =  12'b110000101001;     //233pi/512
   m_cos[233]  =  12'b000100011111;     //233pi/512
   m_sin[234]  =  12'b110000100111;     //234pi/512
   m_cos[234]  =  12'b000100011001;     //234pi/512
   m_sin[235]  =  12'b110000100110;     //235pi/512
   m_cos[235]  =  12'b000100010100;     //235pi/512
   m_sin[236]  =  12'b110000100100;     //236pi/512
   m_cos[236]  =  12'b000100001110;     //236pi/512
   m_sin[237]  =  12'b110000100011;     //237pi/512
   m_cos[237]  =  12'b000100001001;     //237pi/512
   m_sin[238]  =  12'b110000100001;     //238pi/512
   m_cos[238]  =  12'b000100000011;     //238pi/512
   m_sin[239]  =  12'b110000100000;     //239pi/512
   m_cos[239]  =  12'b000011111110;     //239pi/512
   m_sin[240]  =  12'b110000011111;     //240pi/512
   m_cos[240]  =  12'b000011111000;     //240pi/512
   m_sin[241]  =  12'b110000011101;     //241pi/512
   m_cos[241]  =  12'b000011110011;     //241pi/512
   m_sin[242]  =  12'b110000011100;     //242pi/512
   m_cos[242]  =  12'b000011101101;     //242pi/512
   m_sin[243]  =  12'b110000011011;     //243pi/512
   m_cos[243]  =  12'b000011101000;     //243pi/512
   m_sin[244]  =  12'b110000011001;     //244pi/512
   m_cos[244]  =  12'b000011100010;     //244pi/512
   m_sin[245]  =  12'b110000011000;     //245pi/512
   m_cos[245]  =  12'b000011011101;     //245pi/512
   m_sin[246]  =  12'b110000010111;     //246pi/512
   m_cos[246]  =  12'b000011010111;     //246pi/512
   m_sin[247]  =  12'b110000010110;     //247pi/512
   m_cos[247]  =  12'b000011010010;     //247pi/512
   m_sin[248]  =  12'b110000010101;     //248pi/512
   m_cos[248]  =  12'b000011001100;     //248pi/512
   m_sin[249]  =  12'b110000010100;     //249pi/512
   m_cos[249]  =  12'b000011000111;     //249pi/512
   m_sin[250]  =  12'b110000010010;     //250pi/512
   m_cos[250]  =  12'b000011000001;     //250pi/512
   m_sin[251]  =  12'b110000010001;     //251pi/512
   m_cos[251]  =  12'b000010111100;     //251pi/512
   m_sin[252]  =  12'b110000010000;     //252pi/512
   m_cos[252]  =  12'b000010110110;     //252pi/512
   m_sin[253]  =  12'b110000001111;     //253pi/512
   m_cos[253]  =  12'b000010110000;     //253pi/512
   m_sin[254]  =  12'b110000001110;     //254pi/512
   m_cos[254]  =  12'b000010101011;     //254pi/512
   m_sin[255]  =  12'b110000001110;     //255pi/512
   m_cos[255]  =  12'b000010100101;     //255pi/512
   m_sin[256]  =  12'b110000001101;     //256pi/512
   m_cos[256]  =  12'b000010100000;     //256pi/512
   m_sin[257]  =  12'b110000001100;     //257pi/512
   m_cos[257]  =  12'b000010011010;     //257pi/512
   m_sin[258]  =  12'b110000001011;     //258pi/512
   m_cos[258]  =  12'b000010010101;     //258pi/512
   m_sin[259]  =  12'b110000001010;     //259pi/512
   m_cos[259]  =  12'b000010001111;     //259pi/512
   m_sin[260]  =  12'b110000001001;     //260pi/512
   m_cos[260]  =  12'b000010001001;     //260pi/512
   m_sin[261]  =  12'b110000001001;     //261pi/512
   m_cos[261]  =  12'b000010000100;     //261pi/512
   m_sin[262]  =  12'b110000001000;     //262pi/512
   m_cos[262]  =  12'b000001111110;     //262pi/512
   m_sin[263]  =  12'b110000000111;     //263pi/512
   m_cos[263]  =  12'b000001111000;     //263pi/512
   m_sin[264]  =  12'b110000000111;     //264pi/512
   m_cos[264]  =  12'b000001110011;     //264pi/512
   m_sin[265]  =  12'b110000000110;     //265pi/512
   m_cos[265]  =  12'b000001101101;     //265pi/512
   m_sin[266]  =  12'b110000000101;     //266pi/512
   m_cos[266]  =  12'b000001101000;     //266pi/512
   m_sin[267]  =  12'b110000000101;     //267pi/512
   m_cos[267]  =  12'b000001100010;     //267pi/512
   m_sin[268]  =  12'b110000000100;     //268pi/512
   m_cos[268]  =  12'b000001011100;     //268pi/512
   m_sin[269]  =  12'b110000000100;     //269pi/512
   m_cos[269]  =  12'b000001010111;     //269pi/512
   m_sin[270]  =  12'b110000000011;     //270pi/512
   m_cos[270]  =  12'b000001010001;     //270pi/512
   m_sin[271]  =  12'b110000000011;     //271pi/512
   m_cos[271]  =  12'b000001001011;     //271pi/512
   m_sin[272]  =  12'b110000000010;     //272pi/512
   m_cos[272]  =  12'b000001000110;     //272pi/512
   m_sin[273]  =  12'b110000000010;     //273pi/512
   m_cos[273]  =  12'b000001000000;     //273pi/512
   m_sin[274]  =  12'b110000000010;     //274pi/512
   m_cos[274]  =  12'b000000111011;     //274pi/512
   m_sin[275]  =  12'b110000000001;     //275pi/512
   m_cos[275]  =  12'b000000110101;     //275pi/512
   m_sin[276]  =  12'b110000000001;     //276pi/512
   m_cos[276]  =  12'b000000101111;     //276pi/512
   m_sin[277]  =  12'b110000000001;     //277pi/512
   m_cos[277]  =  12'b000000101010;     //277pi/512
   m_sin[278]  =  12'b110000000001;     //278pi/512
   m_cos[278]  =  12'b000000100100;     //278pi/512
   m_sin[279]  =  12'b110000000000;     //279pi/512
   m_cos[279]  =  12'b000000011110;     //279pi/512
   m_sin[280]  =  12'b110000000000;     //280pi/512
   m_cos[280]  =  12'b000000011001;     //280pi/512
   m_sin[281]  =  12'b110000000000;     //281pi/512
   m_cos[281]  =  12'b000000010011;     //281pi/512
   m_sin[282]  =  12'b110000000000;     //282pi/512
   m_cos[282]  =  12'b000000001101;     //282pi/512
   m_sin[283]  =  12'b110000000000;     //283pi/512
   m_cos[283]  =  12'b000000001000;     //283pi/512
   m_sin[284]  =  12'b110000000000;     //284pi/512
   m_cos[284]  =  12'b000000000010;     //284pi/512
   m_sin[285]  =  12'b110000000000;     //285pi/512
   m_cos[285]  =  12'b111111111101;     //285pi/512
   m_sin[286]  =  12'b110000000000;     //286pi/512
   m_cos[286]  =  12'b111111110111;     //286pi/512
   m_sin[287]  =  12'b110000000000;     //287pi/512
   m_cos[287]  =  12'b111111110010;     //287pi/512
   m_sin[288]  =  12'b110000000000;     //288pi/512
   m_cos[288]  =  12'b111111101100;     //288pi/512
   m_sin[289]  =  12'b110000000000;     //289pi/512
   m_cos[289]  =  12'b111111100110;     //289pi/512
   m_sin[290]  =  12'b110000000000;     //290pi/512
   m_cos[290]  =  12'b111111100001;     //290pi/512
   m_sin[291]  =  12'b110000000001;     //291pi/512
   m_cos[291]  =  12'b111111011011;     //291pi/512
   m_sin[292]  =  12'b110000000001;     //292pi/512
   m_cos[292]  =  12'b111111010101;     //292pi/512
   m_sin[293]  =  12'b110000000001;     //293pi/512
   m_cos[293]  =  12'b111111010000;     //293pi/512
   m_sin[294]  =  12'b110000000001;     //294pi/512
   m_cos[294]  =  12'b111111001010;     //294pi/512
   m_sin[295]  =  12'b110000000010;     //295pi/512
   m_cos[295]  =  12'b111111000100;     //295pi/512
   m_sin[296]  =  12'b110000000010;     //296pi/512
   m_cos[296]  =  12'b111110111111;     //296pi/512
   m_sin[297]  =  12'b110000000010;     //297pi/512
   m_cos[297]  =  12'b111110111001;     //297pi/512
   m_sin[298]  =  12'b110000000011;     //298pi/512
   m_cos[298]  =  12'b111110110011;     //298pi/512
   m_sin[299]  =  12'b110000000011;     //299pi/512
   m_cos[299]  =  12'b111110101110;     //299pi/512
   m_sin[300]  =  12'b110000000100;     //300pi/512
   m_cos[300]  =  12'b111110101000;     //300pi/512
   m_sin[301]  =  12'b110000000100;     //301pi/512
   m_cos[301]  =  12'b111110100011;     //301pi/512
   m_sin[302]  =  12'b110000000101;     //302pi/512
   m_cos[302]  =  12'b111110011101;     //302pi/512
   m_sin[303]  =  12'b110000000101;     //303pi/512
   m_cos[303]  =  12'b111110010111;     //303pi/512
   m_sin[304]  =  12'b110000000110;     //304pi/512
   m_cos[304]  =  12'b111110010010;     //304pi/512
   m_sin[305]  =  12'b110000000111;     //305pi/512
   m_cos[305]  =  12'b111110001100;     //305pi/512
   m_sin[306]  =  12'b110000000111;     //306pi/512
   m_cos[306]  =  12'b111110000110;     //306pi/512
   m_sin[307]  =  12'b110000001000;     //307pi/512
   m_cos[307]  =  12'b111110000001;     //307pi/512
   m_sin[308]  =  12'b110000001001;     //308pi/512
   m_cos[308]  =  12'b111101111011;     //308pi/512
   m_sin[309]  =  12'b110000001001;     //309pi/512
   m_cos[309]  =  12'b111101110110;     //309pi/512
   m_sin[310]  =  12'b110000001010;     //310pi/512
   m_cos[310]  =  12'b111101110000;     //310pi/512
   m_sin[311]  =  12'b110000001011;     //311pi/512
   m_cos[311]  =  12'b111101101010;     //311pi/512
   m_sin[312]  =  12'b110000001100;     //312pi/512
   m_cos[312]  =  12'b111101100101;     //312pi/512
   m_sin[313]  =  12'b110000001101;     //313pi/512
   m_cos[313]  =  12'b111101011111;     //313pi/512
   m_sin[314]  =  12'b110000001110;     //314pi/512
   m_cos[314]  =  12'b111101011010;     //314pi/512
   m_sin[315]  =  12'b110000001111;     //315pi/512
   m_cos[315]  =  12'b111101010100;     //315pi/512
   m_sin[316]  =  12'b110000010000;     //316pi/512
   m_cos[316]  =  12'b111101001110;     //316pi/512
   m_sin[317]  =  12'b110000010001;     //317pi/512
   m_cos[317]  =  12'b111101001001;     //317pi/512
   m_sin[318]  =  12'b110000010010;     //318pi/512
   m_cos[318]  =  12'b111101000011;     //318pi/512
   m_sin[319]  =  12'b110000010011;     //319pi/512
   m_cos[319]  =  12'b111100111110;     //319pi/512
   m_sin[320]  =  12'b110000010100;     //320pi/512
   m_cos[320]  =  12'b111100111000;     //320pi/512
   m_sin[321]  =  12'b110000010101;     //321pi/512
   m_cos[321]  =  12'b111100110011;     //321pi/512
   m_sin[322]  =  12'b110000010110;     //322pi/512
   m_cos[322]  =  12'b111100101101;     //322pi/512
   m_sin[323]  =  12'b110000010111;     //323pi/512
   m_cos[323]  =  12'b111100101000;     //323pi/512
   m_sin[324]  =  12'b110000011000;     //324pi/512
   m_cos[324]  =  12'b111100100010;     //324pi/512
   m_sin[325]  =  12'b110000011010;     //325pi/512
   m_cos[325]  =  12'b111100011101;     //325pi/512
   m_sin[326]  =  12'b110000011011;     //326pi/512
   m_cos[326]  =  12'b111100010111;     //326pi/512
   m_sin[327]  =  12'b110000011100;     //327pi/512
   m_cos[327]  =  12'b111100010010;     //327pi/512
   m_sin[328]  =  12'b110000011101;     //328pi/512
   m_cos[328]  =  12'b111100001100;     //328pi/512
   m_sin[329]  =  12'b110000011111;     //329pi/512
   m_cos[329]  =  12'b111100000111;     //329pi/512
   m_sin[330]  =  12'b110000100000;     //330pi/512
   m_cos[330]  =  12'b111100000001;     //330pi/512
   m_sin[331]  =  12'b110000100010;     //331pi/512
   m_cos[331]  =  12'b111011111100;     //331pi/512
   m_sin[332]  =  12'b110000100011;     //332pi/512
   m_cos[332]  =  12'b111011110110;     //332pi/512
   m_sin[333]  =  12'b110000100101;     //333pi/512
   m_cos[333]  =  12'b111011110001;     //333pi/512
   m_sin[334]  =  12'b110000100110;     //334pi/512
   m_cos[334]  =  12'b111011101011;     //334pi/512
   m_sin[335]  =  12'b110000101000;     //335pi/512
   m_cos[335]  =  12'b111011100110;     //335pi/512
   m_sin[336]  =  12'b110000101001;     //336pi/512
   m_cos[336]  =  12'b111011100000;     //336pi/512
   m_sin[337]  =  12'b110000101011;     //337pi/512
   m_cos[337]  =  12'b111011011011;     //337pi/512
   m_sin[338]  =  12'b110000101100;     //338pi/512
   m_cos[338]  =  12'b111011010110;     //338pi/512
   m_sin[339]  =  12'b110000101110;     //339pi/512
   m_cos[339]  =  12'b111011010000;     //339pi/512
   m_sin[340]  =  12'b110000110000;     //340pi/512
   m_cos[340]  =  12'b111011001011;     //340pi/512
   m_sin[341]  =  12'b110000110010;     //341pi/512
   m_cos[341]  =  12'b111011000101;     //341pi/512
   m_sin[342]  =  12'b110000110011;     //342pi/512
   m_cos[342]  =  12'b111011000000;     //342pi/512
   m_sin[343]  =  12'b110000110101;     //343pi/512
   m_cos[343]  =  12'b111010111011;     //343pi/512
   m_sin[344]  =  12'b110000110111;     //344pi/512
   m_cos[344]  =  12'b111010110101;     //344pi/512
   m_sin[345]  =  12'b110000111001;     //345pi/512
   m_cos[345]  =  12'b111010110000;     //345pi/512
   m_sin[346]  =  12'b110000111011;     //346pi/512
   m_cos[346]  =  12'b111010101011;     //346pi/512
   m_sin[347]  =  12'b110000111100;     //347pi/512
   m_cos[347]  =  12'b111010100101;     //347pi/512
   m_sin[348]  =  12'b110000111110;     //348pi/512
   m_cos[348]  =  12'b111010100000;     //348pi/512
   m_sin[349]  =  12'b110001000000;     //349pi/512
   m_cos[349]  =  12'b111010011011;     //349pi/512
   m_sin[350]  =  12'b110001000010;     //350pi/512
   m_cos[350]  =  12'b111010010101;     //350pi/512
   m_sin[351]  =  12'b110001000100;     //351pi/512
   m_cos[351]  =  12'b111010010000;     //351pi/512
   m_sin[352]  =  12'b110001000110;     //352pi/512
   m_cos[352]  =  12'b111010001011;     //352pi/512
   m_sin[353]  =  12'b110001001001;     //353pi/512
   m_cos[353]  =  12'b111010000110;     //353pi/512
   m_sin[354]  =  12'b110001001011;     //354pi/512
   m_cos[354]  =  12'b111010000000;     //354pi/512
   m_sin[355]  =  12'b110001001101;     //355pi/512
   m_cos[355]  =  12'b111001111011;     //355pi/512
   m_sin[356]  =  12'b110001001111;     //356pi/512
   m_cos[356]  =  12'b111001110110;     //356pi/512
   m_sin[357]  =  12'b110001010001;     //357pi/512
   m_cos[357]  =  12'b111001110001;     //357pi/512
   m_sin[358]  =  12'b110001010011;     //358pi/512
   m_cos[358]  =  12'b111001101011;     //358pi/512
   m_sin[359]  =  12'b110001010110;     //359pi/512
   m_cos[359]  =  12'b111001100110;     //359pi/512
   m_sin[360]  =  12'b110001011000;     //360pi/512
   m_cos[360]  =  12'b111001100001;     //360pi/512
   m_sin[361]  =  12'b110001011010;     //361pi/512
   m_cos[361]  =  12'b111001011100;     //361pi/512
   m_sin[362]  =  12'b110001011100;     //362pi/512
   m_cos[362]  =  12'b111001010111;     //362pi/512
   m_sin[363]  =  12'b110001011111;     //363pi/512
   m_cos[363]  =  12'b111001010010;     //363pi/512
   m_sin[364]  =  12'b110001100001;     //364pi/512
   m_cos[364]  =  12'b111001001100;     //364pi/512
   m_sin[365]  =  12'b110001100100;     //365pi/512
   m_cos[365]  =  12'b111001000111;     //365pi/512
   m_sin[366]  =  12'b110001100110;     //366pi/512
   m_cos[366]  =  12'b111001000010;     //366pi/512
   m_sin[367]  =  12'b110001101001;     //367pi/512
   m_cos[367]  =  12'b111000111101;     //367pi/512
   m_sin[368]  =  12'b110001101011;     //368pi/512
   m_cos[368]  =  12'b111000111000;     //368pi/512
   m_sin[369]  =  12'b110001101110;     //369pi/512
   m_cos[369]  =  12'b111000110011;     //369pi/512
   m_sin[370]  =  12'b110001110000;     //370pi/512
   m_cos[370]  =  12'b111000101110;     //370pi/512
   m_sin[371]  =  12'b110001110011;     //371pi/512
   m_cos[371]  =  12'b111000101001;     //371pi/512
   m_sin[372]  =  12'b110001110101;     //372pi/512
   m_cos[372]  =  12'b111000100100;     //372pi/512
   m_sin[373]  =  12'b110001111000;     //373pi/512
   m_cos[373]  =  12'b111000011111;     //373pi/512
   m_sin[374]  =  12'b110001111011;     //374pi/512
   m_cos[374]  =  12'b111000011010;     //374pi/512
   m_sin[375]  =  12'b110001111101;     //375pi/512
   m_cos[375]  =  12'b111000010101;     //375pi/512
   m_sin[376]  =  12'b110010000000;     //376pi/512
   m_cos[376]  =  12'b111000010000;     //376pi/512
   m_sin[377]  =  12'b110010000011;     //377pi/512
   m_cos[377]  =  12'b111000001011;     //377pi/512
   m_sin[378]  =  12'b110010000110;     //378pi/512
   m_cos[378]  =  12'b111000000110;     //378pi/512
   m_sin[379]  =  12'b110010001000;     //379pi/512
   m_cos[379]  =  12'b111000000001;     //379pi/512
   m_sin[380]  =  12'b110010001011;     //380pi/512
   m_cos[380]  =  12'b110111111100;     //380pi/512
   m_sin[381]  =  12'b110010001110;     //381pi/512
   m_cos[381]  =  12'b110111110111;     //381pi/512
   m_sin[382]  =  12'b110010010001;     //382pi/512
   m_cos[382]  =  12'b110111110011;     //382pi/512
   m_sin[383]  =  12'b110010010100;     //383pi/512
   m_cos[383]  =  12'b110111101110;     //383pi/512
   m_sin[384]  =  12'b110010010111;     //384pi/512
   m_cos[384]  =  12'b110111101001;     //384pi/512
   m_sin[385]  =  12'b110010011010;     //385pi/512
   m_cos[385]  =  12'b110111100100;     //385pi/512
   m_sin[386]  =  12'b110010011101;     //386pi/512
   m_cos[386]  =  12'b110111011111;     //386pi/512
   m_sin[387]  =  12'b110010100000;     //387pi/512
   m_cos[387]  =  12'b110111011011;     //387pi/512
   m_sin[388]  =  12'b110010100011;     //388pi/512
   m_cos[388]  =  12'b110111010110;     //388pi/512
   m_sin[389]  =  12'b110010100110;     //389pi/512
   m_cos[389]  =  12'b110111010001;     //389pi/512
   m_sin[390]  =  12'b110010101001;     //390pi/512
   m_cos[390]  =  12'b110111001100;     //390pi/512
   m_sin[391]  =  12'b110010101100;     //391pi/512
   m_cos[391]  =  12'b110111001000;     //391pi/512
   m_sin[392]  =  12'b110010101111;     //392pi/512
   m_cos[392]  =  12'b110111000011;     //392pi/512
   m_sin[393]  =  12'b110010110011;     //393pi/512
   m_cos[393]  =  12'b110110111110;     //393pi/512
   m_sin[394]  =  12'b110010110110;     //394pi/512
   m_cos[394]  =  12'b110110111010;     //394pi/512
   m_sin[395]  =  12'b110010111001;     //395pi/512
   m_cos[395]  =  12'b110110110101;     //395pi/512
   m_sin[396]  =  12'b110010111100;     //396pi/512
   m_cos[396]  =  12'b110110110000;     //396pi/512
   m_sin[397]  =  12'b110011000000;     //397pi/512
   m_cos[397]  =  12'b110110101100;     //397pi/512
   m_sin[398]  =  12'b110011000011;     //398pi/512
   m_cos[398]  =  12'b110110100111;     //398pi/512
   m_sin[399]  =  12'b110011000110;     //399pi/512
   m_cos[399]  =  12'b110110100011;     //399pi/512
   m_sin[400]  =  12'b110011001010;     //400pi/512
   m_cos[400]  =  12'b110110011110;     //400pi/512
   m_sin[401]  =  12'b110011001101;     //401pi/512
   m_cos[401]  =  12'b110110011001;     //401pi/512
   m_sin[402]  =  12'b110011010000;     //402pi/512
   m_cos[402]  =  12'b110110010101;     //402pi/512
   m_sin[403]  =  12'b110011010100;     //403pi/512
   m_cos[403]  =  12'b110110010000;     //403pi/512
   m_sin[404]  =  12'b110011010111;     //404pi/512
   m_cos[404]  =  12'b110110001100;     //404pi/512
   m_sin[405]  =  12'b110011011011;     //405pi/512
   m_cos[405]  =  12'b110110001000;     //405pi/512
   m_sin[406]  =  12'b110011011110;     //406pi/512
   m_cos[406]  =  12'b110110000011;     //406pi/512
   m_sin[407]  =  12'b110011100010;     //407pi/512
   m_cos[407]  =  12'b110101111111;     //407pi/512
   m_sin[408]  =  12'b110011100101;     //408pi/512
   m_cos[408]  =  12'b110101111010;     //408pi/512
   m_sin[409]  =  12'b110011101001;     //409pi/512
   m_cos[409]  =  12'b110101110110;     //409pi/512
   m_sin[410]  =  12'b110011101100;     //410pi/512
   m_cos[410]  =  12'b110101110010;     //410pi/512
   m_sin[411]  =  12'b110011110000;     //411pi/512
   m_cos[411]  =  12'b110101101101;     //411pi/512
   m_sin[412]  =  12'b110011110100;     //412pi/512
   m_cos[412]  =  12'b110101101001;     //412pi/512
   m_sin[413]  =  12'b110011110111;     //413pi/512
   m_cos[413]  =  12'b110101100101;     //413pi/512
   m_sin[414]  =  12'b110011111011;     //414pi/512
   m_cos[414]  =  12'b110101100000;     //414pi/512
   m_sin[415]  =  12'b110011111111;     //415pi/512
   m_cos[415]  =  12'b110101011100;     //415pi/512
   m_sin[416]  =  12'b110100000011;     //416pi/512
   m_cos[416]  =  12'b110101011000;     //416pi/512
   m_sin[417]  =  12'b110100000110;     //417pi/512
   m_cos[417]  =  12'b110101010100;     //417pi/512
   m_sin[418]  =  12'b110100001010;     //418pi/512
   m_cos[418]  =  12'b110101001111;     //418pi/512
   m_sin[419]  =  12'b110100001110;     //419pi/512
   m_cos[419]  =  12'b110101001011;     //419pi/512
   m_sin[420]  =  12'b110100010010;     //420pi/512
   m_cos[420]  =  12'b110101000111;     //420pi/512
   m_sin[421]  =  12'b110100010110;     //421pi/512
   m_cos[421]  =  12'b110101000011;     //421pi/512
   m_sin[422]  =  12'b110100011010;     //422pi/512
   m_cos[422]  =  12'b110100111111;     //422pi/512
   m_sin[423]  =  12'b110100011101;     //423pi/512
   m_cos[423]  =  12'b110100111011;     //423pi/512
   m_sin[424]  =  12'b110100100001;     //424pi/512
   m_cos[424]  =  12'b110100110111;     //424pi/512
   m_sin[425]  =  12'b110100100101;     //425pi/512
   m_cos[425]  =  12'b110100110011;     //425pi/512
   m_sin[426]  =  12'b110100101001;     //426pi/512
   m_cos[426]  =  12'b110100101111;     //426pi/512
   m_sin[427]  =  12'b110100101101;     //427pi/512
   m_cos[427]  =  12'b110100101011;     //427pi/512
   m_sin[428]  =  12'b110100110001;     //428pi/512
   m_cos[428]  =  12'b110100100111;     //428pi/512
   m_sin[429]  =  12'b110100110101;     //429pi/512
   m_cos[429]  =  12'b110100100011;     //429pi/512
   m_sin[430]  =  12'b110100111001;     //430pi/512
   m_cos[430]  =  12'b110100011111;     //430pi/512
   m_sin[431]  =  12'b110100111101;     //431pi/512
   m_cos[431]  =  12'b110100011011;     //431pi/512
   m_sin[432]  =  12'b110101000010;     //432pi/512
   m_cos[432]  =  12'b110100010111;     //432pi/512
   m_sin[433]  =  12'b110101000110;     //433pi/512
   m_cos[433]  =  12'b110100010011;     //433pi/512
   m_sin[434]  =  12'b110101001010;     //434pi/512
   m_cos[434]  =  12'b110100001111;     //434pi/512
   m_sin[435]  =  12'b110101001110;     //435pi/512
   m_cos[435]  =  12'b110100001011;     //435pi/512
   m_sin[436]  =  12'b110101010010;     //436pi/512
   m_cos[436]  =  12'b110100001000;     //436pi/512
   m_sin[437]  =  12'b110101010110;     //437pi/512
   m_cos[437]  =  12'b110100000100;     //437pi/512
   m_sin[438]  =  12'b110101011011;     //438pi/512
   m_cos[438]  =  12'b110100000000;     //438pi/512
   m_sin[439]  =  12'b110101011111;     //439pi/512
   m_cos[439]  =  12'b110011111100;     //439pi/512
   m_sin[440]  =  12'b110101100011;     //440pi/512
   m_cos[440]  =  12'b110011111001;     //440pi/512
   m_sin[441]  =  12'b110101100111;     //441pi/512
   m_cos[441]  =  12'b110011110101;     //441pi/512
   m_sin[442]  =  12'b110101101100;     //442pi/512
   m_cos[442]  =  12'b110011110001;     //442pi/512
   m_sin[443]  =  12'b110101110000;     //443pi/512
   m_cos[443]  =  12'b110011101110;     //443pi/512
   m_sin[444]  =  12'b110101110100;     //444pi/512
   m_cos[444]  =  12'b110011101010;     //444pi/512
   m_sin[445]  =  12'b110101111001;     //445pi/512
   m_cos[445]  =  12'b110011100110;     //445pi/512
   m_sin[446]  =  12'b110101111101;     //446pi/512
   m_cos[446]  =  12'b110011100011;     //446pi/512
   m_sin[447]  =  12'b110110000010;     //447pi/512
   m_cos[447]  =  12'b110011011111;     //447pi/512
   m_sin[448]  =  12'b110110000110;     //448pi/512
   m_cos[448]  =  12'b110011011100;     //448pi/512
   m_sin[449]  =  12'b110110001010;     //449pi/512
   m_cos[449]  =  12'b110011011000;     //449pi/512
   m_sin[450]  =  12'b110110001111;     //450pi/512
   m_cos[450]  =  12'b110011010101;     //450pi/512
   m_sin[451]  =  12'b110110010011;     //451pi/512
   m_cos[451]  =  12'b110011010001;     //451pi/512
   m_sin[452]  =  12'b110110011000;     //452pi/512
   m_cos[452]  =  12'b110011001110;     //452pi/512
   m_sin[453]  =  12'b110110011100;     //453pi/512
   m_cos[453]  =  12'b110011001011;     //453pi/512
   m_sin[454]  =  12'b110110100001;     //454pi/512
   m_cos[454]  =  12'b110011000111;     //454pi/512
   m_sin[455]  =  12'b110110100110;     //455pi/512
   m_cos[455]  =  12'b110011000100;     //455pi/512
   m_sin[456]  =  12'b110110101010;     //456pi/512
   m_cos[456]  =  12'b110011000001;     //456pi/512
   m_sin[457]  =  12'b110110101111;     //457pi/512
   m_cos[457]  =  12'b110010111101;     //457pi/512
   m_sin[458]  =  12'b110110110011;     //458pi/512
   m_cos[458]  =  12'b110010111010;     //458pi/512
   m_sin[459]  =  12'b110110111000;     //459pi/512
   m_cos[459]  =  12'b110010110111;     //459pi/512
   m_sin[460]  =  12'b110110111101;     //460pi/512
   m_cos[460]  =  12'b110010110100;     //460pi/512
   m_sin[461]  =  12'b110111000001;     //461pi/512
   m_cos[461]  =  12'b110010110000;     //461pi/512
   m_sin[462]  =  12'b110111000110;     //462pi/512
   m_cos[462]  =  12'b110010101101;     //462pi/512
   m_sin[463]  =  12'b110111001011;     //463pi/512
   m_cos[463]  =  12'b110010101010;     //463pi/512
   m_sin[464]  =  12'b110111001111;     //464pi/512
   m_cos[464]  =  12'b110010100111;     //464pi/512
   m_sin[465]  =  12'b110111010100;     //465pi/512
   m_cos[465]  =  12'b110010100100;     //465pi/512
   m_sin[466]  =  12'b110111011001;     //466pi/512
   m_cos[466]  =  12'b110010100001;     //466pi/512
   m_sin[467]  =  12'b110111011110;     //467pi/512
   m_cos[467]  =  12'b110010011110;     //467pi/512
   m_sin[468]  =  12'b110111100011;     //468pi/512
   m_cos[468]  =  12'b110010011011;     //468pi/512
   m_sin[469]  =  12'b110111100111;     //469pi/512
   m_cos[469]  =  12'b110010011000;     //469pi/512
   m_sin[470]  =  12'b110111101100;     //470pi/512
   m_cos[470]  =  12'b110010010101;     //470pi/512
   m_sin[471]  =  12'b110111110001;     //471pi/512
   m_cos[471]  =  12'b110010010010;     //471pi/512
   m_sin[472]  =  12'b110111110110;     //472pi/512
   m_cos[472]  =  12'b110010001111;     //472pi/512
   m_sin[473]  =  12'b110111111011;     //473pi/512
   m_cos[473]  =  12'b110010001100;     //473pi/512
   m_sin[474]  =  12'b111000000000;     //474pi/512
   m_cos[474]  =  12'b110010001001;     //474pi/512
   m_sin[475]  =  12'b111000000101;     //475pi/512
   m_cos[475]  =  12'b110010000111;     //475pi/512
   m_sin[476]  =  12'b111000001001;     //476pi/512
   m_cos[476]  =  12'b110010000100;     //476pi/512
   m_sin[477]  =  12'b111000001110;     //477pi/512
   m_cos[477]  =  12'b110010000001;     //477pi/512
   m_sin[478]  =  12'b111000010011;     //478pi/512
   m_cos[478]  =  12'b110001111110;     //478pi/512
   m_sin[479]  =  12'b111000011000;     //479pi/512
   m_cos[479]  =  12'b110001111100;     //479pi/512
   m_sin[480]  =  12'b111000011101;     //480pi/512
   m_cos[480]  =  12'b110001111001;     //480pi/512
   m_sin[481]  =  12'b111000100010;     //481pi/512
   m_cos[481]  =  12'b110001110110;     //481pi/512
   m_sin[482]  =  12'b111000100111;     //482pi/512
   m_cos[482]  =  12'b110001110100;     //482pi/512
   m_sin[483]  =  12'b111000101100;     //483pi/512
   m_cos[483]  =  12'b110001110001;     //483pi/512
   m_sin[484]  =  12'b111000110001;     //484pi/512
   m_cos[484]  =  12'b110001101110;     //484pi/512
   m_sin[485]  =  12'b111000110110;     //485pi/512
   m_cos[485]  =  12'b110001101100;     //485pi/512
   m_sin[486]  =  12'b111000111011;     //486pi/512
   m_cos[486]  =  12'b110001101001;     //486pi/512
   m_sin[487]  =  12'b111001000001;     //487pi/512
   m_cos[487]  =  12'b110001100111;     //487pi/512
   m_sin[488]  =  12'b111001000110;     //488pi/512
   m_cos[488]  =  12'b110001100100;     //488pi/512
   m_sin[489]  =  12'b111001001011;     //489pi/512
   m_cos[489]  =  12'b110001100010;     //489pi/512
   m_sin[490]  =  12'b111001010000;     //490pi/512
   m_cos[490]  =  12'b110001100000;     //490pi/512
   m_sin[491]  =  12'b111001010101;     //491pi/512
   m_cos[491]  =  12'b110001011101;     //491pi/512
   m_sin[492]  =  12'b111001011010;     //492pi/512
   m_cos[492]  =  12'b110001011011;     //492pi/512
   m_sin[493]  =  12'b111001011111;     //493pi/512
   m_cos[493]  =  12'b110001011001;     //493pi/512
   m_sin[494]  =  12'b111001100100;     //494pi/512
   m_cos[494]  =  12'b110001010110;     //494pi/512
   m_sin[495]  =  12'b111001101010;     //495pi/512
   m_cos[495]  =  12'b110001010100;     //495pi/512
   m_sin[496]  =  12'b111001101111;     //496pi/512
   m_cos[496]  =  12'b110001010010;     //496pi/512
   m_sin[497]  =  12'b111001110100;     //497pi/512
   m_cos[497]  =  12'b110001010000;     //497pi/512
   m_sin[498]  =  12'b111001111001;     //498pi/512
   m_cos[498]  =  12'b110001001101;     //498pi/512
   m_sin[499]  =  12'b111001111111;     //499pi/512
   m_cos[499]  =  12'b110001001011;     //499pi/512
   m_sin[500]  =  12'b111010000100;     //500pi/512
   m_cos[500]  =  12'b110001001001;     //500pi/512
   m_sin[501]  =  12'b111010001001;     //501pi/512
   m_cos[501]  =  12'b110001000111;     //501pi/512
   m_sin[502]  =  12'b111010001110;     //502pi/512
   m_cos[502]  =  12'b110001000101;     //502pi/512
   m_sin[503]  =  12'b111010010100;     //503pi/512
   m_cos[503]  =  12'b110001000011;     //503pi/512
   m_sin[504]  =  12'b111010011001;     //504pi/512
   m_cos[504]  =  12'b110001000001;     //504pi/512
   m_sin[505]  =  12'b111010011110;     //505pi/512
   m_cos[505]  =  12'b110000111111;     //505pi/512
   m_sin[506]  =  12'b111010100011;     //506pi/512
   m_cos[506]  =  12'b110000111101;     //506pi/512
   m_sin[507]  =  12'b111010101001;     //507pi/512
   m_cos[507]  =  12'b110000111011;     //507pi/512
   m_sin[508]  =  12'b111010101110;     //508pi/512
   m_cos[508]  =  12'b110000111001;     //508pi/512
   m_sin[509]  =  12'b111010110011;     //509pi/512
   m_cos[509]  =  12'b110000110111;     //509pi/512
   m_sin[510]  =  12'b111010111001;     //510pi/512
   m_cos[510]  =  12'b110000110110;     //510pi/512
   m_sin[511]  =  12'b111010111110;     //511pi/512
   m_cos[511]  =  12'b110000110100;     //511pi/512
end
endmodule
