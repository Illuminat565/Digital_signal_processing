module  M_TWIDLE_14_bit #(parameter stage_FFT = 2, SIZE =10, word_length_tw = 14) (
    input            clk,
    input            en_rd, 
    input   [stage_FFT-2:0]   rd_ptr_angle,

    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );

reg signed [word_length_tw-1:0]  m_cos  [511:0];
reg signed [word_length_tw-1:0]  m_sin  [511:0];

wire [8:0] rd_ptr  =  rd_ptr_angle << (10-stage_FFT);


//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd ) begin
                  cos_data           <= m_cos   [rd_ptr];
                  sin_data           <= m_sin   [rd_ptr];
             end 
        end
//----------------------------------------------------------------------------------------
initial begin

   m_sin[0]  =  14'b00000000000000;     //0pi/512
   m_cos[0]  =  14'b01000000000000;     //0pi/512
   m_sin[1]  =  14'b11111111101100;     //1pi/512
   m_cos[1]  =  14'b00111111111111;     //1pi/512
   m_sin[2]  =  14'b11111111011000;     //2pi/512
   m_cos[2]  =  14'b00111111111111;     //2pi/512
   m_sin[3]  =  14'b11111111000100;     //3pi/512
   m_cos[3]  =  14'b00111111111111;     //3pi/512
   m_sin[4]  =  14'b11111110110000;     //4pi/512
   m_cos[4]  =  14'b00111111111111;     //4pi/512
   m_sin[5]  =  14'b11111110011011;     //5pi/512
   m_cos[5]  =  14'b00111111111110;     //5pi/512
   m_sin[6]  =  14'b11111110000111;     //6pi/512
   m_cos[6]  =  14'b00111111111110;     //6pi/512
   m_sin[7]  =  14'b11111101110011;     //7pi/512
   m_cos[7]  =  14'b00111111111101;     //7pi/512
   m_sin[8]  =  14'b11111101011111;     //8pi/512
   m_cos[8]  =  14'b00111111111100;     //8pi/512
   m_sin[9]  =  14'b11111101001011;     //9pi/512
   m_cos[9]  =  14'b00111111111100;     //9pi/512
   m_sin[10]  =  14'b11111100110111;     //10pi/512
   m_cos[10]  =  14'b00111111111011;     //10pi/512
   m_sin[11]  =  14'b11111100100011;     //11pi/512
   m_cos[11]  =  14'b00111111111010;     //11pi/512
   m_sin[12]  =  14'b11111100001111;     //12pi/512
   m_cos[12]  =  14'b00111111111000;     //12pi/512
   m_sin[13]  =  14'b11111011111011;     //13pi/512
   m_cos[13]  =  14'b00111111110111;     //13pi/512
   m_sin[14]  =  14'b11111011100111;     //14pi/512
   m_cos[14]  =  14'b00111111110110;     //14pi/512
   m_sin[15]  =  14'b11111011010011;     //15pi/512
   m_cos[15]  =  14'b00111111110100;     //15pi/512
   m_sin[16]  =  14'b11111010111111;     //16pi/512
   m_cos[16]  =  14'b00111111110011;     //16pi/512
   m_sin[17]  =  14'b11111010101011;     //17pi/512
   m_cos[17]  =  14'b00111111110001;     //17pi/512
   m_sin[18]  =  14'b11111010010111;     //18pi/512
   m_cos[18]  =  14'b00111111110000;     //18pi/512
   m_sin[19]  =  14'b11111010000011;     //19pi/512
   m_cos[19]  =  14'b00111111101110;     //19pi/512
   m_sin[20]  =  14'b11111001101111;     //20pi/512
   m_cos[20]  =  14'b00111111101100;     //20pi/512
   m_sin[21]  =  14'b11111001011011;     //21pi/512
   m_cos[21]  =  14'b00111111101010;     //21pi/512
   m_sin[22]  =  14'b11111001000111;     //22pi/512
   m_cos[22]  =  14'b00111111101000;     //22pi/512
   m_sin[23]  =  14'b11111000110011;     //23pi/512
   m_cos[23]  =  14'b00111111100101;     //23pi/512
   m_sin[24]  =  14'b11111000011111;     //24pi/512
   m_cos[24]  =  14'b00111111100011;     //24pi/512
   m_sin[25]  =  14'b11111000001011;     //25pi/512
   m_cos[25]  =  14'b00111111100001;     //25pi/512
   m_sin[26]  =  14'b11110111110111;     //26pi/512
   m_cos[26]  =  14'b00111111011110;     //26pi/512
   m_sin[27]  =  14'b11110111100011;     //27pi/512
   m_cos[27]  =  14'b00111111011100;     //27pi/512
   m_sin[28]  =  14'b11110111001111;     //28pi/512
   m_cos[28]  =  14'b00111111011001;     //28pi/512
   m_sin[29]  =  14'b11110110111011;     //29pi/512
   m_cos[29]  =  14'b00111111010110;     //29pi/512
   m_sin[30]  =  14'b11110110100111;     //30pi/512
   m_cos[30]  =  14'b00111111010011;     //30pi/512
   m_sin[31]  =  14'b11110110010011;     //31pi/512
   m_cos[31]  =  14'b00111111010000;     //31pi/512
   m_sin[32]  =  14'b11110101111111;     //32pi/512
   m_cos[32]  =  14'b00111111001101;     //32pi/512
   m_sin[33]  =  14'b11110101101011;     //33pi/512
   m_cos[33]  =  14'b00111111001010;     //33pi/512
   m_sin[34]  =  14'b11110101011000;     //34pi/512
   m_cos[34]  =  14'b00111111000111;     //34pi/512
   m_sin[35]  =  14'b11110101000100;     //35pi/512
   m_cos[35]  =  14'b00111111000011;     //35pi/512
   m_sin[36]  =  14'b11110100110000;     //36pi/512
   m_cos[36]  =  14'b00111111000000;     //36pi/512
   m_sin[37]  =  14'b11110100011100;     //37pi/512
   m_cos[37]  =  14'b00111110111100;     //37pi/512
   m_sin[38]  =  14'b11110100001000;     //38pi/512
   m_cos[38]  =  14'b00111110111000;     //38pi/512
   m_sin[39]  =  14'b11110011110101;     //39pi/512
   m_cos[39]  =  14'b00111110110101;     //39pi/512
   m_sin[40]  =  14'b11110011100001;     //40pi/512
   m_cos[40]  =  14'b00111110110001;     //40pi/512
   m_sin[41]  =  14'b11110011001101;     //41pi/512
   m_cos[41]  =  14'b00111110101101;     //41pi/512
   m_sin[42]  =  14'b11110010111010;     //42pi/512
   m_cos[42]  =  14'b00111110101001;     //42pi/512
   m_sin[43]  =  14'b11110010100110;     //43pi/512
   m_cos[43]  =  14'b00111110100101;     //43pi/512
   m_sin[44]  =  14'b11110010010010;     //44pi/512
   m_cos[44]  =  14'b00111110100000;     //44pi/512
   m_sin[45]  =  14'b11110001111111;     //45pi/512
   m_cos[45]  =  14'b00111110011100;     //45pi/512
   m_sin[46]  =  14'b11110001101011;     //46pi/512
   m_cos[46]  =  14'b00111110011000;     //46pi/512
   m_sin[47]  =  14'b11110001010111;     //47pi/512
   m_cos[47]  =  14'b00111110010011;     //47pi/512
   m_sin[48]  =  14'b11110001000100;     //48pi/512
   m_cos[48]  =  14'b00111110001110;     //48pi/512
   m_sin[49]  =  14'b11110000110000;     //49pi/512
   m_cos[49]  =  14'b00111110001010;     //49pi/512
   m_sin[50]  =  14'b11110000011101;     //50pi/512
   m_cos[50]  =  14'b00111110000101;     //50pi/512
   m_sin[51]  =  14'b11110000001001;     //51pi/512
   m_cos[51]  =  14'b00111110000000;     //51pi/512
   m_sin[52]  =  14'b11101111110110;     //52pi/512
   m_cos[52]  =  14'b00111101111011;     //52pi/512
   m_sin[53]  =  14'b11101111100010;     //53pi/512
   m_cos[53]  =  14'b00111101110110;     //53pi/512
   m_sin[54]  =  14'b11101111001111;     //54pi/512
   m_cos[54]  =  14'b00111101110000;     //54pi/512
   m_sin[55]  =  14'b11101110111100;     //55pi/512
   m_cos[55]  =  14'b00111101101011;     //55pi/512
   m_sin[56]  =  14'b11101110101000;     //56pi/512
   m_cos[56]  =  14'b00111101100110;     //56pi/512
   m_sin[57]  =  14'b11101110010101;     //57pi/512
   m_cos[57]  =  14'b00111101100000;     //57pi/512
   m_sin[58]  =  14'b11101110000010;     //58pi/512
   m_cos[58]  =  14'b00111101011011;     //58pi/512
   m_sin[59]  =  14'b11101101101110;     //59pi/512
   m_cos[59]  =  14'b00111101010101;     //59pi/512
   m_sin[60]  =  14'b11101101011011;     //60pi/512
   m_cos[60]  =  14'b00111101001111;     //60pi/512
   m_sin[61]  =  14'b11101101001000;     //61pi/512
   m_cos[61]  =  14'b00111101001001;     //61pi/512
   m_sin[62]  =  14'b11101100110101;     //62pi/512
   m_cos[62]  =  14'b00111101000011;     //62pi/512
   m_sin[63]  =  14'b11101100100001;     //63pi/512
   m_cos[63]  =  14'b00111100111101;     //63pi/512
   m_sin[64]  =  14'b11101100001110;     //64pi/512
   m_cos[64]  =  14'b00111100110111;     //64pi/512
   m_sin[65]  =  14'b11101011111011;     //65pi/512
   m_cos[65]  =  14'b00111100110001;     //65pi/512
   m_sin[66]  =  14'b11101011101000;     //66pi/512
   m_cos[66]  =  14'b00111100101010;     //66pi/512
   m_sin[67]  =  14'b11101011010101;     //67pi/512
   m_cos[67]  =  14'b00111100100100;     //67pi/512
   m_sin[68]  =  14'b11101011000010;     //68pi/512
   m_cos[68]  =  14'b00111100011101;     //68pi/512
   m_sin[69]  =  14'b11101010101111;     //69pi/512
   m_cos[69]  =  14'b00111100010111;     //69pi/512
   m_sin[70]  =  14'b11101010011100;     //70pi/512
   m_cos[70]  =  14'b00111100010000;     //70pi/512
   m_sin[71]  =  14'b11101010001001;     //71pi/512
   m_cos[71]  =  14'b00111100001001;     //71pi/512
   m_sin[72]  =  14'b11101001110110;     //72pi/512
   m_cos[72]  =  14'b00111100000010;     //72pi/512
   m_sin[73]  =  14'b11101001100011;     //73pi/512
   m_cos[73]  =  14'b00111011111011;     //73pi/512
   m_sin[74]  =  14'b11101001010001;     //74pi/512
   m_cos[74]  =  14'b00111011110100;     //74pi/512
   m_sin[75]  =  14'b11101000111110;     //75pi/512
   m_cos[75]  =  14'b00111011101101;     //75pi/512
   m_sin[76]  =  14'b11101000101011;     //76pi/512
   m_cos[76]  =  14'b00111011100110;     //76pi/512
   m_sin[77]  =  14'b11101000011000;     //77pi/512
   m_cos[77]  =  14'b00111011011110;     //77pi/512
   m_sin[78]  =  14'b11101000000110;     //78pi/512
   m_cos[78]  =  14'b00111011010111;     //78pi/512
   m_sin[79]  =  14'b11100111110011;     //79pi/512
   m_cos[79]  =  14'b00111011001111;     //79pi/512
   m_sin[80]  =  14'b11100111100001;     //80pi/512
   m_cos[80]  =  14'b00111011001000;     //80pi/512
   m_sin[81]  =  14'b11100111001110;     //81pi/512
   m_cos[81]  =  14'b00111011000000;     //81pi/512
   m_sin[82]  =  14'b11100110111011;     //82pi/512
   m_cos[82]  =  14'b00111010111000;     //82pi/512
   m_sin[83]  =  14'b11100110101001;     //83pi/512
   m_cos[83]  =  14'b00111010110000;     //83pi/512
   m_sin[84]  =  14'b11100110010111;     //84pi/512
   m_cos[84]  =  14'b00111010101000;     //84pi/512
   m_sin[85]  =  14'b11100110000100;     //85pi/512
   m_cos[85]  =  14'b00111010100000;     //85pi/512
   m_sin[86]  =  14'b11100101110010;     //86pi/512
   m_cos[86]  =  14'b00111010011000;     //86pi/512
   m_sin[87]  =  14'b11100101011111;     //87pi/512
   m_cos[87]  =  14'b00111010010000;     //87pi/512
   m_sin[88]  =  14'b11100101001101;     //88pi/512
   m_cos[88]  =  14'b00111010000111;     //88pi/512
   m_sin[89]  =  14'b11100100111011;     //89pi/512
   m_cos[89]  =  14'b00111001111111;     //89pi/512
   m_sin[90]  =  14'b11100100101001;     //90pi/512
   m_cos[90]  =  14'b00111001110110;     //90pi/512
   m_sin[91]  =  14'b11100100010111;     //91pi/512
   m_cos[91]  =  14'b00111001101110;     //91pi/512
   m_sin[92]  =  14'b11100100000100;     //92pi/512
   m_cos[92]  =  14'b00111001100101;     //92pi/512
   m_sin[93]  =  14'b11100011110010;     //93pi/512
   m_cos[93]  =  14'b00111001011100;     //93pi/512
   m_sin[94]  =  14'b11100011100000;     //94pi/512
   m_cos[94]  =  14'b00111001010011;     //94pi/512
   m_sin[95]  =  14'b11100011001110;     //95pi/512
   m_cos[95]  =  14'b00111001001010;     //95pi/512
   m_sin[96]  =  14'b11100010111100;     //96pi/512
   m_cos[96]  =  14'b00111001000001;     //96pi/512
   m_sin[97]  =  14'b11100010101011;     //97pi/512
   m_cos[97]  =  14'b00111000111000;     //97pi/512
   m_sin[98]  =  14'b11100010011001;     //98pi/512
   m_cos[98]  =  14'b00111000101111;     //98pi/512
   m_sin[99]  =  14'b11100010000111;     //99pi/512
   m_cos[99]  =  14'b00111000100101;     //99pi/512
   m_sin[100]  =  14'b11100001110101;     //100pi/512
   m_cos[100]  =  14'b00111000011100;     //100pi/512
   m_sin[101]  =  14'b11100001100011;     //101pi/512
   m_cos[101]  =  14'b00111000010010;     //101pi/512
   m_sin[102]  =  14'b11100001010010;     //102pi/512
   m_cos[102]  =  14'b00111000001001;     //102pi/512
   m_sin[103]  =  14'b11100001000000;     //103pi/512
   m_cos[103]  =  14'b00110111111111;     //103pi/512
   m_sin[104]  =  14'b11100000101111;     //104pi/512
   m_cos[104]  =  14'b00110111110101;     //104pi/512
   m_sin[105]  =  14'b11100000011101;     //105pi/512
   m_cos[105]  =  14'b00110111101011;     //105pi/512
   m_sin[106]  =  14'b11100000001100;     //106pi/512
   m_cos[106]  =  14'b00110111100001;     //106pi/512
   m_sin[107]  =  14'b11011111111010;     //107pi/512
   m_cos[107]  =  14'b00110111010111;     //107pi/512
   m_sin[108]  =  14'b11011111101001;     //108pi/512
   m_cos[108]  =  14'b00110111001101;     //108pi/512
   m_sin[109]  =  14'b11011111011000;     //109pi/512
   m_cos[109]  =  14'b00110111000011;     //109pi/512
   m_sin[110]  =  14'b11011111000110;     //110pi/512
   m_cos[110]  =  14'b00110110111001;     //110pi/512
   m_sin[111]  =  14'b11011110110101;     //111pi/512
   m_cos[111]  =  14'b00110110101110;     //111pi/512
   m_sin[112]  =  14'b11011110100100;     //112pi/512
   m_cos[112]  =  14'b00110110100100;     //112pi/512
   m_sin[113]  =  14'b11011110010011;     //113pi/512
   m_cos[113]  =  14'b00110110011001;     //113pi/512
   m_sin[114]  =  14'b11011110000010;     //114pi/512
   m_cos[114]  =  14'b00110110001111;     //114pi/512
   m_sin[115]  =  14'b11011101110001;     //115pi/512
   m_cos[115]  =  14'b00110110000100;     //115pi/512
   m_sin[116]  =  14'b11011101100000;     //116pi/512
   m_cos[116]  =  14'b00110101111001;     //116pi/512
   m_sin[117]  =  14'b11011101001111;     //117pi/512
   m_cos[117]  =  14'b00110101101110;     //117pi/512
   m_sin[118]  =  14'b11011100111110;     //118pi/512
   m_cos[118]  =  14'b00110101100011;     //118pi/512
   m_sin[119]  =  14'b11011100101101;     //119pi/512
   m_cos[119]  =  14'b00110101011000;     //119pi/512
   m_sin[120]  =  14'b11011100011100;     //120pi/512
   m_cos[120]  =  14'b00110101001101;     //120pi/512
   m_sin[121]  =  14'b11011100001100;     //121pi/512
   m_cos[121]  =  14'b00110101000010;     //121pi/512
   m_sin[122]  =  14'b11011011111011;     //122pi/512
   m_cos[122]  =  14'b00110100110111;     //122pi/512
   m_sin[123]  =  14'b11011011101010;     //123pi/512
   m_cos[123]  =  14'b00110100101011;     //123pi/512
   m_sin[124]  =  14'b11011011011010;     //124pi/512
   m_cos[124]  =  14'b00110100100000;     //124pi/512
   m_sin[125]  =  14'b11011011001001;     //125pi/512
   m_cos[125]  =  14'b00110100010100;     //125pi/512
   m_sin[126]  =  14'b11011010111001;     //126pi/512
   m_cos[126]  =  14'b00110100001001;     //126pi/512
   m_sin[127]  =  14'b11011010101001;     //127pi/512
   m_cos[127]  =  14'b00110011111101;     //127pi/512
   m_sin[128]  =  14'b11011010011000;     //128pi/512
   m_cos[128]  =  14'b00110011110001;     //128pi/512
   m_sin[129]  =  14'b11011010001000;     //129pi/512
   m_cos[129]  =  14'b00110011100101;     //129pi/512
   m_sin[130]  =  14'b11011001111000;     //130pi/512
   m_cos[130]  =  14'b00110011011001;     //130pi/512
   m_sin[131]  =  14'b11011001101000;     //131pi/512
   m_cos[131]  =  14'b00110011001101;     //131pi/512
   m_sin[132]  =  14'b11011001011000;     //132pi/512
   m_cos[132]  =  14'b00110011000001;     //132pi/512
   m_sin[133]  =  14'b11011001001000;     //133pi/512
   m_cos[133]  =  14'b00110010110101;     //133pi/512
   m_sin[134]  =  14'b11011000111000;     //134pi/512
   m_cos[134]  =  14'b00110010101001;     //134pi/512
   m_sin[135]  =  14'b11011000101000;     //135pi/512
   m_cos[135]  =  14'b00110010011101;     //135pi/512
   m_sin[136]  =  14'b11011000011000;     //136pi/512
   m_cos[136]  =  14'b00110010010000;     //136pi/512
   m_sin[137]  =  14'b11011000001000;     //137pi/512
   m_cos[137]  =  14'b00110010000100;     //137pi/512
   m_sin[138]  =  14'b11010111111001;     //138pi/512
   m_cos[138]  =  14'b00110001110111;     //138pi/512
   m_sin[139]  =  14'b11010111101001;     //139pi/512
   m_cos[139]  =  14'b00110001101010;     //139pi/512
   m_sin[140]  =  14'b11010111011010;     //140pi/512
   m_cos[140]  =  14'b00110001011110;     //140pi/512
   m_sin[141]  =  14'b11010111001010;     //141pi/512
   m_cos[141]  =  14'b00110001010001;     //141pi/512
   m_sin[142]  =  14'b11010110111011;     //142pi/512
   m_cos[142]  =  14'b00110001000100;     //142pi/512
   m_sin[143]  =  14'b11010110101011;     //143pi/512
   m_cos[143]  =  14'b00110000110111;     //143pi/512
   m_sin[144]  =  14'b11010110011100;     //144pi/512
   m_cos[144]  =  14'b00110000101010;     //144pi/512
   m_sin[145]  =  14'b11010110001101;     //145pi/512
   m_cos[145]  =  14'b00110000011101;     //145pi/512
   m_sin[146]  =  14'b11010101111101;     //146pi/512
   m_cos[146]  =  14'b00110000010000;     //146pi/512
   m_sin[147]  =  14'b11010101101110;     //147pi/512
   m_cos[147]  =  14'b00110000000011;     //147pi/512
   m_sin[148]  =  14'b11010101011111;     //148pi/512
   m_cos[148]  =  14'b00101111110101;     //148pi/512
   m_sin[149]  =  14'b11010101010000;     //149pi/512
   m_cos[149]  =  14'b00101111101000;     //149pi/512
   m_sin[150]  =  14'b11010101000001;     //150pi/512
   m_cos[150]  =  14'b00101111011010;     //150pi/512
   m_sin[151]  =  14'b11010100110010;     //151pi/512
   m_cos[151]  =  14'b00101111001101;     //151pi/512
   m_sin[152]  =  14'b11010100100100;     //152pi/512
   m_cos[152]  =  14'b00101110111111;     //152pi/512
   m_sin[153]  =  14'b11010100010101;     //153pi/512
   m_cos[153]  =  14'b00101110110010;     //153pi/512
   m_sin[154]  =  14'b11010100000110;     //154pi/512
   m_cos[154]  =  14'b00101110100100;     //154pi/512
   m_sin[155]  =  14'b11010011111000;     //155pi/512
   m_cos[155]  =  14'b00101110010110;     //155pi/512
   m_sin[156]  =  14'b11010011101001;     //156pi/512
   m_cos[156]  =  14'b00101110001000;     //156pi/512
   m_sin[157]  =  14'b11010011011011;     //157pi/512
   m_cos[157]  =  14'b00101101111010;     //157pi/512
   m_sin[158]  =  14'b11010011001100;     //158pi/512
   m_cos[158]  =  14'b00101101101100;     //158pi/512
   m_sin[159]  =  14'b11010010111110;     //159pi/512
   m_cos[159]  =  14'b00101101011110;     //159pi/512
   m_sin[160]  =  14'b11010010110000;     //160pi/512
   m_cos[160]  =  14'b00101101010000;     //160pi/512
   m_sin[161]  =  14'b11010010100010;     //161pi/512
   m_cos[161]  =  14'b00101101000010;     //161pi/512
   m_sin[162]  =  14'b11010010010011;     //162pi/512
   m_cos[162]  =  14'b00101100110011;     //162pi/512
   m_sin[163]  =  14'b11010010000101;     //163pi/512
   m_cos[163]  =  14'b00101100100101;     //163pi/512
   m_sin[164]  =  14'b11010001110111;     //164pi/512
   m_cos[164]  =  14'b00101100010110;     //164pi/512
   m_sin[165]  =  14'b11010001101001;     //165pi/512
   m_cos[165]  =  14'b00101100001000;     //165pi/512
   m_sin[166]  =  14'b11010001011100;     //166pi/512
   m_cos[166]  =  14'b00101011111001;     //166pi/512
   m_sin[167]  =  14'b11010001001110;     //167pi/512
   m_cos[167]  =  14'b00101011101011;     //167pi/512
   m_sin[168]  =  14'b11010001000000;     //168pi/512
   m_cos[168]  =  14'b00101011011100;     //168pi/512
   m_sin[169]  =  14'b11010000110011;     //169pi/512
   m_cos[169]  =  14'b00101011001101;     //169pi/512
   m_sin[170]  =  14'b11010000100101;     //170pi/512
   m_cos[170]  =  14'b00101010111110;     //170pi/512
   m_sin[171]  =  14'b11010000011000;     //171pi/512
   m_cos[171]  =  14'b00101010101111;     //171pi/512
   m_sin[172]  =  14'b11010000001010;     //172pi/512
   m_cos[172]  =  14'b00101010100000;     //172pi/512
   m_sin[173]  =  14'b11001111111101;     //173pi/512
   m_cos[173]  =  14'b00101010010001;     //173pi/512
   m_sin[174]  =  14'b11001111110000;     //174pi/512
   m_cos[174]  =  14'b00101010000010;     //174pi/512
   m_sin[175]  =  14'b11001111100010;     //175pi/512
   m_cos[175]  =  14'b00101001110011;     //175pi/512
   m_sin[176]  =  14'b11001111010101;     //176pi/512
   m_cos[176]  =  14'b00101001100100;     //176pi/512
   m_sin[177]  =  14'b11001111001000;     //177pi/512
   m_cos[177]  =  14'b00101001010100;     //177pi/512
   m_sin[178]  =  14'b11001110111011;     //178pi/512
   m_cos[178]  =  14'b00101001000101;     //178pi/512
   m_sin[179]  =  14'b11001110101111;     //179pi/512
   m_cos[179]  =  14'b00101000110101;     //179pi/512
   m_sin[180]  =  14'b11001110100010;     //180pi/512
   m_cos[180]  =  14'b00101000100110;     //180pi/512
   m_sin[181]  =  14'b11001110010101;     //181pi/512
   m_cos[181]  =  14'b00101000010110;     //181pi/512
   m_sin[182]  =  14'b11001110001000;     //182pi/512
   m_cos[182]  =  14'b00101000000111;     //182pi/512
   m_sin[183]  =  14'b11001101111100;     //183pi/512
   m_cos[183]  =  14'b00100111110111;     //183pi/512
   m_sin[184]  =  14'b11001101101111;     //184pi/512
   m_cos[184]  =  14'b00100111100111;     //184pi/512
   m_sin[185]  =  14'b11001101100011;     //185pi/512
   m_cos[185]  =  14'b00100111010111;     //185pi/512
   m_sin[186]  =  14'b11001101010111;     //186pi/512
   m_cos[186]  =  14'b00100111001000;     //186pi/512
   m_sin[187]  =  14'b11001101001010;     //187pi/512
   m_cos[187]  =  14'b00100110111000;     //187pi/512
   m_sin[188]  =  14'b11001100111110;     //188pi/512
   m_cos[188]  =  14'b00100110101000;     //188pi/512
   m_sin[189]  =  14'b11001100110010;     //189pi/512
   m_cos[189]  =  14'b00100110011000;     //189pi/512
   m_sin[190]  =  14'b11001100100110;     //190pi/512
   m_cos[190]  =  14'b00100110000111;     //190pi/512
   m_sin[191]  =  14'b11001100011010;     //191pi/512
   m_cos[191]  =  14'b00100101110111;     //191pi/512
   m_sin[192]  =  14'b11001100001110;     //192pi/512
   m_cos[192]  =  14'b00100101100111;     //192pi/512
   m_sin[193]  =  14'b11001100000010;     //193pi/512
   m_cos[193]  =  14'b00100101010111;     //193pi/512
   m_sin[194]  =  14'b11001011110111;     //194pi/512
   m_cos[194]  =  14'b00100101000110;     //194pi/512
   m_sin[195]  =  14'b11001011101011;     //195pi/512
   m_cos[195]  =  14'b00100100110110;     //195pi/512
   m_sin[196]  =  14'b11001011100000;     //196pi/512
   m_cos[196]  =  14'b00100100100110;     //196pi/512
   m_sin[197]  =  14'b11001011010100;     //197pi/512
   m_cos[197]  =  14'b00100100010101;     //197pi/512
   m_sin[198]  =  14'b11001011001001;     //198pi/512
   m_cos[198]  =  14'b00100100000100;     //198pi/512
   m_sin[199]  =  14'b11001010111110;     //199pi/512
   m_cos[199]  =  14'b00100011110100;     //199pi/512
   m_sin[200]  =  14'b11001010110010;     //200pi/512
   m_cos[200]  =  14'b00100011100011;     //200pi/512
   m_sin[201]  =  14'b11001010100111;     //201pi/512
   m_cos[201]  =  14'b00100011010010;     //201pi/512
   m_sin[202]  =  14'b11001010011100;     //202pi/512
   m_cos[202]  =  14'b00100011000010;     //202pi/512
   m_sin[203]  =  14'b11001010010001;     //203pi/512
   m_cos[203]  =  14'b00100010110001;     //203pi/512
   m_sin[204]  =  14'b11001010000110;     //204pi/512
   m_cos[204]  =  14'b00100010100000;     //204pi/512
   m_sin[205]  =  14'b11001001111011;     //205pi/512
   m_cos[205]  =  14'b00100010001111;     //205pi/512
   m_sin[206]  =  14'b11001001110001;     //206pi/512
   m_cos[206]  =  14'b00100001111110;     //206pi/512
   m_sin[207]  =  14'b11001001100110;     //207pi/512
   m_cos[207]  =  14'b00100001101101;     //207pi/512
   m_sin[208]  =  14'b11001001011100;     //208pi/512
   m_cos[208]  =  14'b00100001011100;     //208pi/512
   m_sin[209]  =  14'b11001001010001;     //209pi/512
   m_cos[209]  =  14'b00100001001010;     //209pi/512
   m_sin[210]  =  14'b11001001000111;     //210pi/512
   m_cos[210]  =  14'b00100000111001;     //210pi/512
   m_sin[211]  =  14'b11001000111100;     //211pi/512
   m_cos[211]  =  14'b00100000101000;     //211pi/512
   m_sin[212]  =  14'b11001000110010;     //212pi/512
   m_cos[212]  =  14'b00100000010111;     //212pi/512
   m_sin[213]  =  14'b11001000101000;     //213pi/512
   m_cos[213]  =  14'b00100000000101;     //213pi/512
   m_sin[214]  =  14'b11001000011110;     //214pi/512
   m_cos[214]  =  14'b00011111110100;     //214pi/512
   m_sin[215]  =  14'b11001000010100;     //215pi/512
   m_cos[215]  =  14'b00011111100010;     //215pi/512
   m_sin[216]  =  14'b11001000001010;     //216pi/512
   m_cos[216]  =  14'b00011111010001;     //216pi/512
   m_sin[217]  =  14'b11001000000000;     //217pi/512
   m_cos[217]  =  14'b00011110111111;     //217pi/512
   m_sin[218]  =  14'b11000111110111;     //218pi/512
   m_cos[218]  =  14'b00011110101110;     //218pi/512
   m_sin[219]  =  14'b11000111101101;     //219pi/512
   m_cos[219]  =  14'b00011110011100;     //219pi/512
   m_sin[220]  =  14'b11000111100100;     //220pi/512
   m_cos[220]  =  14'b00011110001010;     //220pi/512
   m_sin[221]  =  14'b11000111011010;     //221pi/512
   m_cos[221]  =  14'b00011101111001;     //221pi/512
   m_sin[222]  =  14'b11000111010001;     //222pi/512
   m_cos[222]  =  14'b00011101100111;     //222pi/512
   m_sin[223]  =  14'b11000111001000;     //223pi/512
   m_cos[223]  =  14'b00011101010101;     //223pi/512
   m_sin[224]  =  14'b11000110111110;     //224pi/512
   m_cos[224]  =  14'b00011101000011;     //224pi/512
   m_sin[225]  =  14'b11000110110101;     //225pi/512
   m_cos[225]  =  14'b00011100110001;     //225pi/512
   m_sin[226]  =  14'b11000110101100;     //226pi/512
   m_cos[226]  =  14'b00011100011111;     //226pi/512
   m_sin[227]  =  14'b11000110100011;     //227pi/512
   m_cos[227]  =  14'b00011100001101;     //227pi/512
   m_sin[228]  =  14'b11000110011011;     //228pi/512
   m_cos[228]  =  14'b00011011111011;     //228pi/512
   m_sin[229]  =  14'b11000110010010;     //229pi/512
   m_cos[229]  =  14'b00011011101001;     //229pi/512
   m_sin[230]  =  14'b11000110001001;     //230pi/512
   m_cos[230]  =  14'b00011011010111;     //230pi/512
   m_sin[231]  =  14'b11000110000001;     //231pi/512
   m_cos[231]  =  14'b00011011000101;     //231pi/512
   m_sin[232]  =  14'b11000101111000;     //232pi/512
   m_cos[232]  =  14'b00011010110010;     //232pi/512
   m_sin[233]  =  14'b11000101110000;     //233pi/512
   m_cos[233]  =  14'b00011010100000;     //233pi/512
   m_sin[234]  =  14'b11000101101000;     //234pi/512
   m_cos[234]  =  14'b00011010001110;     //234pi/512
   m_sin[235]  =  14'b11000101011111;     //235pi/512
   m_cos[235]  =  14'b00011001111011;     //235pi/512
   m_sin[236]  =  14'b11000101010111;     //236pi/512
   m_cos[236]  =  14'b00011001101001;     //236pi/512
   m_sin[237]  =  14'b11000101001111;     //237pi/512
   m_cos[237]  =  14'b00011001010111;     //237pi/512
   m_sin[238]  =  14'b11000101000111;     //238pi/512
   m_cos[238]  =  14'b00011001000100;     //238pi/512
   m_sin[239]  =  14'b11000101000000;     //239pi/512
   m_cos[239]  =  14'b00011000110010;     //239pi/512
   m_sin[240]  =  14'b11000100111000;     //240pi/512
   m_cos[240]  =  14'b00011000011111;     //240pi/512
   m_sin[241]  =  14'b11000100110000;     //241pi/512
   m_cos[241]  =  14'b00011000001100;     //241pi/512
   m_sin[242]  =  14'b11000100101001;     //242pi/512
   m_cos[242]  =  14'b00010111111010;     //242pi/512
   m_sin[243]  =  14'b11000100100001;     //243pi/512
   m_cos[243]  =  14'b00010111100111;     //243pi/512
   m_sin[244]  =  14'b11000100011010;     //244pi/512
   m_cos[244]  =  14'b00010111010100;     //244pi/512
   m_sin[245]  =  14'b11000100010010;     //245pi/512
   m_cos[245]  =  14'b00010111000010;     //245pi/512
   m_sin[246]  =  14'b11000100001011;     //246pi/512
   m_cos[246]  =  14'b00010110101111;     //246pi/512
   m_sin[247]  =  14'b11000100000100;     //247pi/512
   m_cos[247]  =  14'b00010110011100;     //247pi/512
   m_sin[248]  =  14'b11000011111101;     //248pi/512
   m_cos[248]  =  14'b00010110001001;     //248pi/512
   m_sin[249]  =  14'b11000011110110;     //249pi/512
   m_cos[249]  =  14'b00010101110110;     //249pi/512
   m_sin[250]  =  14'b11000011101111;     //250pi/512
   m_cos[250]  =  14'b00010101100011;     //250pi/512
   m_sin[251]  =  14'b11000011101001;     //251pi/512
   m_cos[251]  =  14'b00010101010000;     //251pi/512
   m_sin[252]  =  14'b11000011100010;     //252pi/512
   m_cos[252]  =  14'b00010100111101;     //252pi/512
   m_sin[253]  =  14'b11000011011100;     //253pi/512
   m_cos[253]  =  14'b00010100101010;     //253pi/512
   m_sin[254]  =  14'b11000011010101;     //254pi/512
   m_cos[254]  =  14'b00010100010111;     //254pi/512
   m_sin[255]  =  14'b11000011001111;     //255pi/512
   m_cos[255]  =  14'b00010100000100;     //255pi/512
   m_sin[256]  =  14'b11000011001000;     //256pi/512
   m_cos[256]  =  14'b00010011110001;     //256pi/512
   m_sin[257]  =  14'b11000011000010;     //257pi/512
   m_cos[257]  =  14'b00010011011110;     //257pi/512
   m_sin[258]  =  14'b11000010111100;     //258pi/512
   m_cos[258]  =  14'b00010011001011;     //258pi/512
   m_sin[259]  =  14'b11000010110110;     //259pi/512
   m_cos[259]  =  14'b00010010111000;     //259pi/512
   m_sin[260]  =  14'b11000010110000;     //260pi/512
   m_cos[260]  =  14'b00010010100101;     //260pi/512
   m_sin[261]  =  14'b11000010101011;     //261pi/512
   m_cos[261]  =  14'b00010010010001;     //261pi/512
   m_sin[262]  =  14'b11000010100101;     //262pi/512
   m_cos[262]  =  14'b00010001111110;     //262pi/512
   m_sin[263]  =  14'b11000010011111;     //263pi/512
   m_cos[263]  =  14'b00010001101011;     //263pi/512
   m_sin[264]  =  14'b11000010011010;     //264pi/512
   m_cos[264]  =  14'b00010001010111;     //264pi/512
   m_sin[265]  =  14'b11000010010100;     //265pi/512
   m_cos[265]  =  14'b00010001000100;     //265pi/512
   m_sin[266]  =  14'b11000010001111;     //266pi/512
   m_cos[266]  =  14'b00010000110001;     //266pi/512
   m_sin[267]  =  14'b11000010001010;     //267pi/512
   m_cos[267]  =  14'b00010000011101;     //267pi/512
   m_sin[268]  =  14'b11000010000101;     //268pi/512
   m_cos[268]  =  14'b00010000001010;     //268pi/512
   m_sin[269]  =  14'b11000010000000;     //269pi/512
   m_cos[269]  =  14'b00001111110110;     //269pi/512
   m_sin[270]  =  14'b11000001111011;     //270pi/512
   m_cos[270]  =  14'b00001111100011;     //270pi/512
   m_sin[271]  =  14'b11000001110110;     //271pi/512
   m_cos[271]  =  14'b00001111001111;     //271pi/512
   m_sin[272]  =  14'b11000001110001;     //272pi/512
   m_cos[272]  =  14'b00001110111100;     //272pi/512
   m_sin[273]  =  14'b11000001101101;     //273pi/512
   m_cos[273]  =  14'b00001110101000;     //273pi/512
   m_sin[274]  =  14'b11000001101000;     //274pi/512
   m_cos[274]  =  14'b00001110010101;     //274pi/512
   m_sin[275]  =  14'b11000001100100;     //275pi/512
   m_cos[275]  =  14'b00001110000001;     //275pi/512
   m_sin[276]  =  14'b11000001011111;     //276pi/512
   m_cos[276]  =  14'b00001101101101;     //276pi/512
   m_sin[277]  =  14'b11000001011011;     //277pi/512
   m_cos[277]  =  14'b00001101011010;     //277pi/512
   m_sin[278]  =  14'b11000001010111;     //278pi/512
   m_cos[278]  =  14'b00001101000110;     //278pi/512
   m_sin[279]  =  14'b11000001010011;     //279pi/512
   m_cos[279]  =  14'b00001100110010;     //279pi/512
   m_sin[280]  =  14'b11000001001111;     //280pi/512
   m_cos[280]  =  14'b00001100011111;     //280pi/512
   m_sin[281]  =  14'b11000001001011;     //281pi/512
   m_cos[281]  =  14'b00001100001011;     //281pi/512
   m_sin[282]  =  14'b11000001000111;     //282pi/512
   m_cos[282]  =  14'b00001011110111;     //282pi/512
   m_sin[283]  =  14'b11000001000011;     //283pi/512
   m_cos[283]  =  14'b00001011100011;     //283pi/512
   m_sin[284]  =  14'b11000001000000;     //284pi/512
   m_cos[284]  =  14'b00001011010000;     //284pi/512
   m_sin[285]  =  14'b11000000111100;     //285pi/512
   m_cos[285]  =  14'b00001010111100;     //285pi/512
   m_sin[286]  =  14'b11000000111001;     //286pi/512
   m_cos[286]  =  14'b00001010101000;     //286pi/512
   m_sin[287]  =  14'b11000000110110;     //287pi/512
   m_cos[287]  =  14'b00001010010100;     //287pi/512
   m_sin[288]  =  14'b11000000110010;     //288pi/512
   m_cos[288]  =  14'b00001010000000;     //288pi/512
   m_sin[289]  =  14'b11000000101111;     //289pi/512
   m_cos[289]  =  14'b00001001101100;     //289pi/512
   m_sin[290]  =  14'b11000000101100;     //290pi/512
   m_cos[290]  =  14'b00001001011001;     //290pi/512
   m_sin[291]  =  14'b11000000101001;     //291pi/512
   m_cos[291]  =  14'b00001001000101;     //291pi/512
   m_sin[292]  =  14'b11000000100111;     //292pi/512
   m_cos[292]  =  14'b00001000110001;     //292pi/512
   m_sin[293]  =  14'b11000000100100;     //293pi/512
   m_cos[293]  =  14'b00001000011101;     //293pi/512
   m_sin[294]  =  14'b11000000100001;     //294pi/512
   m_cos[294]  =  14'b00001000001001;     //294pi/512
   m_sin[295]  =  14'b11000000011111;     //295pi/512
   m_cos[295]  =  14'b00000111110101;     //295pi/512
   m_sin[296]  =  14'b11000000011100;     //296pi/512
   m_cos[296]  =  14'b00000111100001;     //296pi/512
   m_sin[297]  =  14'b11000000011010;     //297pi/512
   m_cos[297]  =  14'b00000111001101;     //297pi/512
   m_sin[298]  =  14'b11000000011000;     //298pi/512
   m_cos[298]  =  14'b00000110111001;     //298pi/512
   m_sin[299]  =  14'b11000000010110;     //299pi/512
   m_cos[299]  =  14'b00000110100101;     //299pi/512
   m_sin[300]  =  14'b11000000010100;     //300pi/512
   m_cos[300]  =  14'b00000110010001;     //300pi/512
   m_sin[301]  =  14'b11000000010010;     //301pi/512
   m_cos[301]  =  14'b00000101111101;     //301pi/512
   m_sin[302]  =  14'b11000000010000;     //302pi/512
   m_cos[302]  =  14'b00000101101001;     //302pi/512
   m_sin[303]  =  14'b11000000001110;     //303pi/512
   m_cos[303]  =  14'b00000101010101;     //303pi/512
   m_sin[304]  =  14'b11000000001101;     //304pi/512
   m_cos[304]  =  14'b00000101000001;     //304pi/512
   m_sin[305]  =  14'b11000000001011;     //305pi/512
   m_cos[305]  =  14'b00000100101101;     //305pi/512
   m_sin[306]  =  14'b11000000001010;     //306pi/512
   m_cos[306]  =  14'b00000100011001;     //306pi/512
   m_sin[307]  =  14'b11000000001000;     //307pi/512
   m_cos[307]  =  14'b00000100000101;     //307pi/512
   m_sin[308]  =  14'b11000000000111;     //308pi/512
   m_cos[308]  =  14'b00000011110001;     //308pi/512
   m_sin[309]  =  14'b11000000000110;     //309pi/512
   m_cos[309]  =  14'b00000011011101;     //309pi/512
   m_sin[310]  =  14'b11000000000101;     //310pi/512
   m_cos[310]  =  14'b00000011001000;     //310pi/512
   m_sin[311]  =  14'b11000000000100;     //311pi/512
   m_cos[311]  =  14'b00000010110100;     //311pi/512
   m_sin[312]  =  14'b11000000000011;     //312pi/512
   m_cos[312]  =  14'b00000010100000;     //312pi/512
   m_sin[313]  =  14'b11000000000010;     //313pi/512
   m_cos[313]  =  14'b00000010001100;     //313pi/512
   m_sin[314]  =  14'b11000000000010;     //314pi/512
   m_cos[314]  =  14'b00000001111000;     //314pi/512
   m_sin[315]  =  14'b11000000000001;     //315pi/512
   m_cos[315]  =  14'b00000001100100;     //315pi/512
   m_sin[316]  =  14'b11000000000001;     //316pi/512
   m_cos[316]  =  14'b00000001010000;     //316pi/512
   m_sin[317]  =  14'b11000000000000;     //317pi/512
   m_cos[317]  =  14'b00000000111100;     //317pi/512
   m_sin[318]  =  14'b11000000000000;     //318pi/512
   m_cos[318]  =  14'b00000000101000;     //318pi/512
   m_sin[319]  =  14'b11000000000000;     //319pi/512
   m_cos[319]  =  14'b00000000010100;     //319pi/512
   m_sin[320]  =  14'b11000000000000;     //320pi/512
   m_cos[320]  =  14'b00000000000000;     //320pi/512
   m_sin[321]  =  14'b11000000000000;     //321pi/512
   m_cos[321]  =  14'b11111111101100;     //321pi/512
   m_sin[322]  =  14'b11000000000000;     //322pi/512
   m_cos[322]  =  14'b11111111011000;     //322pi/512
   m_sin[323]  =  14'b11000000000000;     //323pi/512
   m_cos[323]  =  14'b11111111000100;     //323pi/512
   m_sin[324]  =  14'b11000000000001;     //324pi/512
   m_cos[324]  =  14'b11111110110000;     //324pi/512
   m_sin[325]  =  14'b11000000000001;     //325pi/512
   m_cos[325]  =  14'b11111110011011;     //325pi/512
   m_sin[326]  =  14'b11000000000010;     //326pi/512
   m_cos[326]  =  14'b11111110000111;     //326pi/512
   m_sin[327]  =  14'b11000000000010;     //327pi/512
   m_cos[327]  =  14'b11111101110011;     //327pi/512
   m_sin[328]  =  14'b11000000000011;     //328pi/512
   m_cos[328]  =  14'b11111101011111;     //328pi/512
   m_sin[329]  =  14'b11000000000100;     //329pi/512
   m_cos[329]  =  14'b11111101001011;     //329pi/512
   m_sin[330]  =  14'b11000000000101;     //330pi/512
   m_cos[330]  =  14'b11111100110111;     //330pi/512
   m_sin[331]  =  14'b11000000000110;     //331pi/512
   m_cos[331]  =  14'b11111100100011;     //331pi/512
   m_sin[332]  =  14'b11000000000111;     //332pi/512
   m_cos[332]  =  14'b11111100001111;     //332pi/512
   m_sin[333]  =  14'b11000000001000;     //333pi/512
   m_cos[333]  =  14'b11111011111011;     //333pi/512
   m_sin[334]  =  14'b11000000001010;     //334pi/512
   m_cos[334]  =  14'b11111011100111;     //334pi/512
   m_sin[335]  =  14'b11000000001011;     //335pi/512
   m_cos[335]  =  14'b11111011010011;     //335pi/512
   m_sin[336]  =  14'b11000000001101;     //336pi/512
   m_cos[336]  =  14'b11111010111111;     //336pi/512
   m_sin[337]  =  14'b11000000001110;     //337pi/512
   m_cos[337]  =  14'b11111010101011;     //337pi/512
   m_sin[338]  =  14'b11000000010000;     //338pi/512
   m_cos[338]  =  14'b11111010010111;     //338pi/512
   m_sin[339]  =  14'b11000000010010;     //339pi/512
   m_cos[339]  =  14'b11111010000011;     //339pi/512
   m_sin[340]  =  14'b11000000010100;     //340pi/512
   m_cos[340]  =  14'b11111001101111;     //340pi/512
   m_sin[341]  =  14'b11000000010110;     //341pi/512
   m_cos[341]  =  14'b11111001011011;     //341pi/512
   m_sin[342]  =  14'b11000000011000;     //342pi/512
   m_cos[342]  =  14'b11111001000111;     //342pi/512
   m_sin[343]  =  14'b11000000011010;     //343pi/512
   m_cos[343]  =  14'b11111000110011;     //343pi/512
   m_sin[344]  =  14'b11000000011100;     //344pi/512
   m_cos[344]  =  14'b11111000011111;     //344pi/512
   m_sin[345]  =  14'b11000000011111;     //345pi/512
   m_cos[345]  =  14'b11111000001011;     //345pi/512
   m_sin[346]  =  14'b11000000100001;     //346pi/512
   m_cos[346]  =  14'b11110111110111;     //346pi/512
   m_sin[347]  =  14'b11000000100100;     //347pi/512
   m_cos[347]  =  14'b11110111100011;     //347pi/512
   m_sin[348]  =  14'b11000000100111;     //348pi/512
   m_cos[348]  =  14'b11110111001111;     //348pi/512
   m_sin[349]  =  14'b11000000101001;     //349pi/512
   m_cos[349]  =  14'b11110110111011;     //349pi/512
   m_sin[350]  =  14'b11000000101100;     //350pi/512
   m_cos[350]  =  14'b11110110100111;     //350pi/512
   m_sin[351]  =  14'b11000000101111;     //351pi/512
   m_cos[351]  =  14'b11110110010011;     //351pi/512
   m_sin[352]  =  14'b11000000110010;     //352pi/512
   m_cos[352]  =  14'b11110101111111;     //352pi/512
   m_sin[353]  =  14'b11000000110110;     //353pi/512
   m_cos[353]  =  14'b11110101101011;     //353pi/512
   m_sin[354]  =  14'b11000000111001;     //354pi/512
   m_cos[354]  =  14'b11110101011000;     //354pi/512
   m_sin[355]  =  14'b11000000111100;     //355pi/512
   m_cos[355]  =  14'b11110101000100;     //355pi/512
   m_sin[356]  =  14'b11000001000000;     //356pi/512
   m_cos[356]  =  14'b11110100110000;     //356pi/512
   m_sin[357]  =  14'b11000001000011;     //357pi/512
   m_cos[357]  =  14'b11110100011100;     //357pi/512
   m_sin[358]  =  14'b11000001000111;     //358pi/512
   m_cos[358]  =  14'b11110100001000;     //358pi/512
   m_sin[359]  =  14'b11000001001011;     //359pi/512
   m_cos[359]  =  14'b11110011110101;     //359pi/512
   m_sin[360]  =  14'b11000001001111;     //360pi/512
   m_cos[360]  =  14'b11110011100001;     //360pi/512
   m_sin[361]  =  14'b11000001010011;     //361pi/512
   m_cos[361]  =  14'b11110011001101;     //361pi/512
   m_sin[362]  =  14'b11000001010111;     //362pi/512
   m_cos[362]  =  14'b11110010111010;     //362pi/512
   m_sin[363]  =  14'b11000001011011;     //363pi/512
   m_cos[363]  =  14'b11110010100110;     //363pi/512
   m_sin[364]  =  14'b11000001011111;     //364pi/512
   m_cos[364]  =  14'b11110010010010;     //364pi/512
   m_sin[365]  =  14'b11000001100100;     //365pi/512
   m_cos[365]  =  14'b11110001111111;     //365pi/512
   m_sin[366]  =  14'b11000001101000;     //366pi/512
   m_cos[366]  =  14'b11110001101011;     //366pi/512
   m_sin[367]  =  14'b11000001101101;     //367pi/512
   m_cos[367]  =  14'b11110001010111;     //367pi/512
   m_sin[368]  =  14'b11000001110001;     //368pi/512
   m_cos[368]  =  14'b11110001000100;     //368pi/512
   m_sin[369]  =  14'b11000001110110;     //369pi/512
   m_cos[369]  =  14'b11110000110000;     //369pi/512
   m_sin[370]  =  14'b11000001111011;     //370pi/512
   m_cos[370]  =  14'b11110000011101;     //370pi/512
   m_sin[371]  =  14'b11000010000000;     //371pi/512
   m_cos[371]  =  14'b11110000001001;     //371pi/512
   m_sin[372]  =  14'b11000010000101;     //372pi/512
   m_cos[372]  =  14'b11101111110110;     //372pi/512
   m_sin[373]  =  14'b11000010001010;     //373pi/512
   m_cos[373]  =  14'b11101111100010;     //373pi/512
   m_sin[374]  =  14'b11000010001111;     //374pi/512
   m_cos[374]  =  14'b11101111001111;     //374pi/512
   m_sin[375]  =  14'b11000010010100;     //375pi/512
   m_cos[375]  =  14'b11101110111100;     //375pi/512
   m_sin[376]  =  14'b11000010011010;     //376pi/512
   m_cos[376]  =  14'b11101110101000;     //376pi/512
   m_sin[377]  =  14'b11000010011111;     //377pi/512
   m_cos[377]  =  14'b11101110010101;     //377pi/512
   m_sin[378]  =  14'b11000010100101;     //378pi/512
   m_cos[378]  =  14'b11101110000010;     //378pi/512
   m_sin[379]  =  14'b11000010101011;     //379pi/512
   m_cos[379]  =  14'b11101101101110;     //379pi/512
   m_sin[380]  =  14'b11000010110000;     //380pi/512
   m_cos[380]  =  14'b11101101011011;     //380pi/512
   m_sin[381]  =  14'b11000010110110;     //381pi/512
   m_cos[381]  =  14'b11101101001000;     //381pi/512
   m_sin[382]  =  14'b11000010111100;     //382pi/512
   m_cos[382]  =  14'b11101100110101;     //382pi/512
   m_sin[383]  =  14'b11000011000010;     //383pi/512
   m_cos[383]  =  14'b11101100100001;     //383pi/512
   m_sin[384]  =  14'b11000011001000;     //384pi/512
   m_cos[384]  =  14'b11101100001110;     //384pi/512
   m_sin[385]  =  14'b11000011001111;     //385pi/512
   m_cos[385]  =  14'b11101011111011;     //385pi/512
   m_sin[386]  =  14'b11000011010101;     //386pi/512
   m_cos[386]  =  14'b11101011101000;     //386pi/512
   m_sin[387]  =  14'b11000011011100;     //387pi/512
   m_cos[387]  =  14'b11101011010101;     //387pi/512
   m_sin[388]  =  14'b11000011100010;     //388pi/512
   m_cos[388]  =  14'b11101011000010;     //388pi/512
   m_sin[389]  =  14'b11000011101001;     //389pi/512
   m_cos[389]  =  14'b11101010101111;     //389pi/512
   m_sin[390]  =  14'b11000011101111;     //390pi/512
   m_cos[390]  =  14'b11101010011100;     //390pi/512
   m_sin[391]  =  14'b11000011110110;     //391pi/512
   m_cos[391]  =  14'b11101010001001;     //391pi/512
   m_sin[392]  =  14'b11000011111101;     //392pi/512
   m_cos[392]  =  14'b11101001110110;     //392pi/512
   m_sin[393]  =  14'b11000100000100;     //393pi/512
   m_cos[393]  =  14'b11101001100011;     //393pi/512
   m_sin[394]  =  14'b11000100001011;     //394pi/512
   m_cos[394]  =  14'b11101001010001;     //394pi/512
   m_sin[395]  =  14'b11000100010010;     //395pi/512
   m_cos[395]  =  14'b11101000111110;     //395pi/512
   m_sin[396]  =  14'b11000100011010;     //396pi/512
   m_cos[396]  =  14'b11101000101011;     //396pi/512
   m_sin[397]  =  14'b11000100100001;     //397pi/512
   m_cos[397]  =  14'b11101000011000;     //397pi/512
   m_sin[398]  =  14'b11000100101001;     //398pi/512
   m_cos[398]  =  14'b11101000000110;     //398pi/512
   m_sin[399]  =  14'b11000100110000;     //399pi/512
   m_cos[399]  =  14'b11100111110011;     //399pi/512
   m_sin[400]  =  14'b11000100111000;     //400pi/512
   m_cos[400]  =  14'b11100111100001;     //400pi/512
   m_sin[401]  =  14'b11000101000000;     //401pi/512
   m_cos[401]  =  14'b11100111001110;     //401pi/512
   m_sin[402]  =  14'b11000101000111;     //402pi/512
   m_cos[402]  =  14'b11100110111011;     //402pi/512
   m_sin[403]  =  14'b11000101001111;     //403pi/512
   m_cos[403]  =  14'b11100110101001;     //403pi/512
   m_sin[404]  =  14'b11000101010111;     //404pi/512
   m_cos[404]  =  14'b11100110010111;     //404pi/512
   m_sin[405]  =  14'b11000101011111;     //405pi/512
   m_cos[405]  =  14'b11100110000100;     //405pi/512
   m_sin[406]  =  14'b11000101101000;     //406pi/512
   m_cos[406]  =  14'b11100101110010;     //406pi/512
   m_sin[407]  =  14'b11000101110000;     //407pi/512
   m_cos[407]  =  14'b11100101011111;     //407pi/512
   m_sin[408]  =  14'b11000101111000;     //408pi/512
   m_cos[408]  =  14'b11100101001101;     //408pi/512
   m_sin[409]  =  14'b11000110000001;     //409pi/512
   m_cos[409]  =  14'b11100100111011;     //409pi/512
   m_sin[410]  =  14'b11000110001001;     //410pi/512
   m_cos[410]  =  14'b11100100101001;     //410pi/512
   m_sin[411]  =  14'b11000110010010;     //411pi/512
   m_cos[411]  =  14'b11100100010111;     //411pi/512
   m_sin[412]  =  14'b11000110011011;     //412pi/512
   m_cos[412]  =  14'b11100100000100;     //412pi/512
   m_sin[413]  =  14'b11000110100011;     //413pi/512
   m_cos[413]  =  14'b11100011110010;     //413pi/512
   m_sin[414]  =  14'b11000110101100;     //414pi/512
   m_cos[414]  =  14'b11100011100000;     //414pi/512
   m_sin[415]  =  14'b11000110110101;     //415pi/512
   m_cos[415]  =  14'b11100011001110;     //415pi/512
   m_sin[416]  =  14'b11000110111110;     //416pi/512
   m_cos[416]  =  14'b11100010111100;     //416pi/512
   m_sin[417]  =  14'b11000111001000;     //417pi/512
   m_cos[417]  =  14'b11100010101011;     //417pi/512
   m_sin[418]  =  14'b11000111010001;     //418pi/512
   m_cos[418]  =  14'b11100010011001;     //418pi/512
   m_sin[419]  =  14'b11000111011010;     //419pi/512
   m_cos[419]  =  14'b11100010000111;     //419pi/512
   m_sin[420]  =  14'b11000111100100;     //420pi/512
   m_cos[420]  =  14'b11100001110101;     //420pi/512
   m_sin[421]  =  14'b11000111101101;     //421pi/512
   m_cos[421]  =  14'b11100001100011;     //421pi/512
   m_sin[422]  =  14'b11000111110111;     //422pi/512
   m_cos[422]  =  14'b11100001010010;     //422pi/512
   m_sin[423]  =  14'b11001000000000;     //423pi/512
   m_cos[423]  =  14'b11100001000000;     //423pi/512
   m_sin[424]  =  14'b11001000001010;     //424pi/512
   m_cos[424]  =  14'b11100000101111;     //424pi/512
   m_sin[425]  =  14'b11001000010100;     //425pi/512
   m_cos[425]  =  14'b11100000011101;     //425pi/512
   m_sin[426]  =  14'b11001000011110;     //426pi/512
   m_cos[426]  =  14'b11100000001100;     //426pi/512
   m_sin[427]  =  14'b11001000101000;     //427pi/512
   m_cos[427]  =  14'b11011111111010;     //427pi/512
   m_sin[428]  =  14'b11001000110010;     //428pi/512
   m_cos[428]  =  14'b11011111101001;     //428pi/512
   m_sin[429]  =  14'b11001000111100;     //429pi/512
   m_cos[429]  =  14'b11011111011000;     //429pi/512
   m_sin[430]  =  14'b11001001000111;     //430pi/512
   m_cos[430]  =  14'b11011111000110;     //430pi/512
   m_sin[431]  =  14'b11001001010001;     //431pi/512
   m_cos[431]  =  14'b11011110110101;     //431pi/512
   m_sin[432]  =  14'b11001001011100;     //432pi/512
   m_cos[432]  =  14'b11011110100100;     //432pi/512
   m_sin[433]  =  14'b11001001100110;     //433pi/512
   m_cos[433]  =  14'b11011110010011;     //433pi/512
   m_sin[434]  =  14'b11001001110001;     //434pi/512
   m_cos[434]  =  14'b11011110000010;     //434pi/512
   m_sin[435]  =  14'b11001001111011;     //435pi/512
   m_cos[435]  =  14'b11011101110001;     //435pi/512
   m_sin[436]  =  14'b11001010000110;     //436pi/512
   m_cos[436]  =  14'b11011101100000;     //436pi/512
   m_sin[437]  =  14'b11001010010001;     //437pi/512
   m_cos[437]  =  14'b11011101001111;     //437pi/512
   m_sin[438]  =  14'b11001010011100;     //438pi/512
   m_cos[438]  =  14'b11011100111110;     //438pi/512
   m_sin[439]  =  14'b11001010100111;     //439pi/512
   m_cos[439]  =  14'b11011100101101;     //439pi/512
   m_sin[440]  =  14'b11001010110010;     //440pi/512
   m_cos[440]  =  14'b11011100011100;     //440pi/512
   m_sin[441]  =  14'b11001010111110;     //441pi/512
   m_cos[441]  =  14'b11011100001100;     //441pi/512
   m_sin[442]  =  14'b11001011001001;     //442pi/512
   m_cos[442]  =  14'b11011011111011;     //442pi/512
   m_sin[443]  =  14'b11001011010100;     //443pi/512
   m_cos[443]  =  14'b11011011101010;     //443pi/512
   m_sin[444]  =  14'b11001011100000;     //444pi/512
   m_cos[444]  =  14'b11011011011010;     //444pi/512
   m_sin[445]  =  14'b11001011101011;     //445pi/512
   m_cos[445]  =  14'b11011011001001;     //445pi/512
   m_sin[446]  =  14'b11001011110111;     //446pi/512
   m_cos[446]  =  14'b11011010111001;     //446pi/512
   m_sin[447]  =  14'b11001100000010;     //447pi/512
   m_cos[447]  =  14'b11011010101001;     //447pi/512
   m_sin[448]  =  14'b11001100001110;     //448pi/512
   m_cos[448]  =  14'b11011010011000;     //448pi/512
   m_sin[449]  =  14'b11001100011010;     //449pi/512
   m_cos[449]  =  14'b11011010001000;     //449pi/512
   m_sin[450]  =  14'b11001100100110;     //450pi/512
   m_cos[450]  =  14'b11011001111000;     //450pi/512
   m_sin[451]  =  14'b11001100110010;     //451pi/512
   m_cos[451]  =  14'b11011001101000;     //451pi/512
   m_sin[452]  =  14'b11001100111110;     //452pi/512
   m_cos[452]  =  14'b11011001011000;     //452pi/512
   m_sin[453]  =  14'b11001101001010;     //453pi/512
   m_cos[453]  =  14'b11011001001000;     //453pi/512
   m_sin[454]  =  14'b11001101010111;     //454pi/512
   m_cos[454]  =  14'b11011000111000;     //454pi/512
   m_sin[455]  =  14'b11001101100011;     //455pi/512
   m_cos[455]  =  14'b11011000101000;     //455pi/512
   m_sin[456]  =  14'b11001101101111;     //456pi/512
   m_cos[456]  =  14'b11011000011000;     //456pi/512
   m_sin[457]  =  14'b11001101111100;     //457pi/512
   m_cos[457]  =  14'b11011000001000;     //457pi/512
   m_sin[458]  =  14'b11001110001000;     //458pi/512
   m_cos[458]  =  14'b11010111111001;     //458pi/512
   m_sin[459]  =  14'b11001110010101;     //459pi/512
   m_cos[459]  =  14'b11010111101001;     //459pi/512
   m_sin[460]  =  14'b11001110100010;     //460pi/512
   m_cos[460]  =  14'b11010111011010;     //460pi/512
   m_sin[461]  =  14'b11001110101111;     //461pi/512
   m_cos[461]  =  14'b11010111001010;     //461pi/512
   m_sin[462]  =  14'b11001110111011;     //462pi/512
   m_cos[462]  =  14'b11010110111011;     //462pi/512
   m_sin[463]  =  14'b11001111001000;     //463pi/512
   m_cos[463]  =  14'b11010110101011;     //463pi/512
   m_sin[464]  =  14'b11001111010101;     //464pi/512
   m_cos[464]  =  14'b11010110011100;     //464pi/512
   m_sin[465]  =  14'b11001111100010;     //465pi/512
   m_cos[465]  =  14'b11010110001101;     //465pi/512
   m_sin[466]  =  14'b11001111110000;     //466pi/512
   m_cos[466]  =  14'b11010101111101;     //466pi/512
   m_sin[467]  =  14'b11001111111101;     //467pi/512
   m_cos[467]  =  14'b11010101101110;     //467pi/512
   m_sin[468]  =  14'b11010000001010;     //468pi/512
   m_cos[468]  =  14'b11010101011111;     //468pi/512
   m_sin[469]  =  14'b11010000011000;     //469pi/512
   m_cos[469]  =  14'b11010101010000;     //469pi/512
   m_sin[470]  =  14'b11010000100101;     //470pi/512
   m_cos[470]  =  14'b11010101000001;     //470pi/512
   m_sin[471]  =  14'b11010000110011;     //471pi/512
   m_cos[471]  =  14'b11010100110010;     //471pi/512
   m_sin[472]  =  14'b11010001000000;     //472pi/512
   m_cos[472]  =  14'b11010100100100;     //472pi/512
   m_sin[473]  =  14'b11010001001110;     //473pi/512
   m_cos[473]  =  14'b11010100010101;     //473pi/512
   m_sin[474]  =  14'b11010001011100;     //474pi/512
   m_cos[474]  =  14'b11010100000110;     //474pi/512
   m_sin[475]  =  14'b11010001101001;     //475pi/512
   m_cos[475]  =  14'b11010011111000;     //475pi/512
   m_sin[476]  =  14'b11010001110111;     //476pi/512
   m_cos[476]  =  14'b11010011101001;     //476pi/512
   m_sin[477]  =  14'b11010010000101;     //477pi/512
   m_cos[477]  =  14'b11010011011011;     //477pi/512
   m_sin[478]  =  14'b11010010010011;     //478pi/512
   m_cos[478]  =  14'b11010011001100;     //478pi/512
   m_sin[479]  =  14'b11010010100010;     //479pi/512
   m_cos[479]  =  14'b11010010111110;     //479pi/512
   m_sin[480]  =  14'b11010010110000;     //480pi/512
   m_cos[480]  =  14'b11010010110000;     //480pi/512
   m_sin[481]  =  14'b11010010111110;     //481pi/512
   m_cos[481]  =  14'b11010010100010;     //481pi/512
   m_sin[482]  =  14'b11010011001100;     //482pi/512
   m_cos[482]  =  14'b11010010010011;     //482pi/512
   m_sin[483]  =  14'b11010011011011;     //483pi/512
   m_cos[483]  =  14'b11010010000101;     //483pi/512
   m_sin[484]  =  14'b11010011101001;     //484pi/512
   m_cos[484]  =  14'b11010001110111;     //484pi/512
   m_sin[485]  =  14'b11010011111000;     //485pi/512
   m_cos[485]  =  14'b11010001101001;     //485pi/512
   m_sin[486]  =  14'b11010100000110;     //486pi/512
   m_cos[486]  =  14'b11010001011100;     //486pi/512
   m_sin[487]  =  14'b11010100010101;     //487pi/512
   m_cos[487]  =  14'b11010001001110;     //487pi/512
   m_sin[488]  =  14'b11010100100100;     //488pi/512
   m_cos[488]  =  14'b11010001000000;     //488pi/512
   m_sin[489]  =  14'b11010100110010;     //489pi/512
   m_cos[489]  =  14'b11010000110011;     //489pi/512
   m_sin[490]  =  14'b11010101000001;     //490pi/512
   m_cos[490]  =  14'b11010000100101;     //490pi/512
   m_sin[491]  =  14'b11010101010000;     //491pi/512
   m_cos[491]  =  14'b11010000011000;     //491pi/512
   m_sin[492]  =  14'b11010101011111;     //492pi/512
   m_cos[492]  =  14'b11010000001010;     //492pi/512
   m_sin[493]  =  14'b11010101101110;     //493pi/512
   m_cos[493]  =  14'b11001111111101;     //493pi/512
   m_sin[494]  =  14'b11010101111101;     //494pi/512
   m_cos[494]  =  14'b11001111110000;     //494pi/512
   m_sin[495]  =  14'b11010110001101;     //495pi/512
   m_cos[495]  =  14'b11001111100010;     //495pi/512
   m_sin[496]  =  14'b11010110011100;     //496pi/512
   m_cos[496]  =  14'b11001111010101;     //496pi/512
   m_sin[497]  =  14'b11010110101011;     //497pi/512
   m_cos[497]  =  14'b11001111001000;     //497pi/512
   m_sin[498]  =  14'b11010110111011;     //498pi/512
   m_cos[498]  =  14'b11001110111011;     //498pi/512
   m_sin[499]  =  14'b11010111001010;     //499pi/512
   m_cos[499]  =  14'b11001110101111;     //499pi/512
   m_sin[500]  =  14'b11010111011010;     //500pi/512
   m_cos[500]  =  14'b11001110100010;     //500pi/512
   m_sin[501]  =  14'b11010111101001;     //501pi/512
   m_cos[501]  =  14'b11001110010101;     //501pi/512
   m_sin[502]  =  14'b11010111111001;     //502pi/512
   m_cos[502]  =  14'b11001110001000;     //502pi/512
   m_sin[503]  =  14'b11011000001000;     //503pi/512
   m_cos[503]  =  14'b11001101111100;     //503pi/512
   m_sin[504]  =  14'b11011000011000;     //504pi/512
   m_cos[504]  =  14'b11001101101111;     //504pi/512
   m_sin[505]  =  14'b11011000101000;     //505pi/512
   m_cos[505]  =  14'b11001101100011;     //505pi/512
   m_sin[506]  =  14'b11011000111000;     //506pi/512
   m_cos[506]  =  14'b11001101010111;     //506pi/512
   m_sin[507]  =  14'b11011001001000;     //507pi/512
   m_cos[507]  =  14'b11001101001010;     //507pi/512
   m_sin[508]  =  14'b11011001011000;     //508pi/512
   m_cos[508]  =  14'b11001100111110;     //508pi/512
   m_sin[509]  =  14'b11011001101000;     //509pi/512
   m_cos[509]  =  14'b11001100110010;     //509pi/512
   m_sin[510]  =  14'b11011001111000;     //510pi/512
   m_cos[510]  =  14'b11001100100110;     //510pi/512
   m_sin[511]  =  14'b11011010001000;     //511pi/512
   m_cos[511]  =  14'b11001100011010;     //511pi/512
end
endmodule