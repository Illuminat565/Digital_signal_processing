module  TWIDLE_8_bit  (
    input   [10:0]   rd_ptr_angle,

    output  signed [7:0]   cos_data,
    output  signed [7:0]   sin_data
 );

wire signed [7:0]  cos  [511:0];
wire signed [7:0]  sin  [511:0];

assign cos_data =    cos [rd_ptr_angle];
assign sin_data =    sin [rd_ptr_angle];

   assign sin[0]  =  8'b00000000;     //0pi/512
  assign cos[0]  =  8'b01000000;     //0pi/512
  assign sin[1]  =  8'b00000000;     //1pi/512
  assign cos[1]  =  8'b00111111;     //1pi/512
  assign sin[2]  =  8'b11111111;     //2pi/512
  assign cos[2]  =  8'b00111111;     //2pi/512
  assign sin[3]  =  8'b11111111;     //3pi/512
  assign cos[3]  =  8'b00111111;     //3pi/512
  assign sin[4]  =  8'b11111110;     //4pi/512
  assign cos[4]  =  8'b00111111;     //4pi/512
  assign sin[5]  =  8'b11111110;     //5pi/512
  assign cos[5]  =  8'b00111111;     //5pi/512
  assign sin[6]  =  8'b11111110;     //6pi/512
  assign cos[6]  =  8'b00111111;     //6pi/512
  assign sin[7]  =  8'b11111101;     //7pi/512
  assign cos[7]  =  8'b00111111;     //7pi/512
  assign sin[8]  =  8'b11111101;     //8pi/512
  assign cos[8]  =  8'b00111111;     //8pi/512
  assign sin[9]  =  8'b11111100;     //9pi/512
  assign cos[9]  =  8'b00111111;     //9pi/512
  assign sin[10]  =  8'b11111100;     //10pi/512
  assign cos[10]  =  8'b00111111;     //10pi/512
  assign sin[11]  =  8'b11111100;     //11pi/512
  assign cos[11]  =  8'b00111111;     //11pi/512
  assign sin[12]  =  8'b11111011;     //12pi/512
  assign cos[12]  =  8'b00111111;     //12pi/512
  assign sin[13]  =  8'b11111011;     //13pi/512
  assign cos[13]  =  8'b00111111;     //13pi/512
  assign sin[14]  =  8'b11111011;     //14pi/512
  assign cos[14]  =  8'b00111111;     //14pi/512
  assign sin[15]  =  8'b11111010;     //15pi/512
  assign cos[15]  =  8'b00111111;     //15pi/512
  assign sin[16]  =  8'b11111010;     //16pi/512
  assign cos[16]  =  8'b00111111;     //16pi/512
  assign sin[17]  =  8'b11111001;     //17pi/512
  assign cos[17]  =  8'b00111111;     //17pi/512
  assign sin[18]  =  8'b11111001;     //18pi/512
  assign cos[18]  =  8'b00111111;     //18pi/512
  assign sin[19]  =  8'b11111001;     //19pi/512
  assign cos[19]  =  8'b00111111;     //19pi/512
  assign sin[20]  =  8'b11111000;     //20pi/512
  assign cos[20]  =  8'b00111111;     //20pi/512
  assign sin[21]  =  8'b11111000;     //21pi/512
  assign cos[21]  =  8'b00111111;     //21pi/512
  assign sin[22]  =  8'b11110111;     //22pi/512
  assign cos[22]  =  8'b00111111;     //22pi/512
  assign sin[23]  =  8'b11110111;     //23pi/512
  assign cos[23]  =  8'b00111111;     //23pi/512
  assign sin[24]  =  8'b11110111;     //24pi/512
  assign cos[24]  =  8'b00111111;     //24pi/512
  assign sin[25]  =  8'b11110110;     //25pi/512
  assign cos[25]  =  8'b00111111;     //25pi/512
  assign sin[26]  =  8'b11110110;     //26pi/512
  assign cos[26]  =  8'b00111111;     //26pi/512
  assign sin[27]  =  8'b11110101;     //27pi/512
  assign cos[27]  =  8'b00111111;     //27pi/512
  assign sin[28]  =  8'b11110101;     //28pi/512
  assign cos[28]  =  8'b00111111;     //28pi/512
  assign sin[29]  =  8'b11110101;     //29pi/512
  assign cos[29]  =  8'b00111110;     //29pi/512
  assign sin[30]  =  8'b11110100;     //30pi/512
  assign cos[30]  =  8'b00111110;     //30pi/512
  assign sin[31]  =  8'b11110100;     //31pi/512
  assign cos[31]  =  8'b00111110;     //31pi/512
  assign sin[32]  =  8'b11110100;     //32pi/512
  assign cos[32]  =  8'b00111110;     //32pi/512
  assign sin[33]  =  8'b11110011;     //33pi/512
  assign cos[33]  =  8'b00111110;     //33pi/512
  assign sin[34]  =  8'b11110011;     //34pi/512
  assign cos[34]  =  8'b00111110;     //34pi/512
  assign sin[35]  =  8'b11110010;     //35pi/512
  assign cos[35]  =  8'b00111110;     //35pi/512
  assign sin[36]  =  8'b11110010;     //36pi/512
  assign cos[36]  =  8'b00111110;     //36pi/512
  assign sin[37]  =  8'b11110010;     //37pi/512
  assign cos[37]  =  8'b00111110;     //37pi/512
  assign sin[38]  =  8'b11110001;     //38pi/512
  assign cos[38]  =  8'b00111110;     //38pi/512
  assign sin[39]  =  8'b11110001;     //39pi/512
  assign cos[39]  =  8'b00111110;     //39pi/512
  assign sin[40]  =  8'b11110000;     //40pi/512
  assign cos[40]  =  8'b00111110;     //40pi/512
  assign sin[41]  =  8'b11110000;     //41pi/512
  assign cos[41]  =  8'b00111101;     //41pi/512
  assign sin[42]  =  8'b11110000;     //42pi/512
  assign cos[42]  =  8'b00111101;     //42pi/512
  assign sin[43]  =  8'b11101111;     //43pi/512
  assign cos[43]  =  8'b00111101;     //43pi/512
  assign sin[44]  =  8'b11101111;     //44pi/512
  assign cos[44]  =  8'b00111101;     //44pi/512
  assign sin[45]  =  8'b11101111;     //45pi/512
  assign cos[45]  =  8'b00111101;     //45pi/512
  assign sin[46]  =  8'b11101110;     //46pi/512
  assign cos[46]  =  8'b00111101;     //46pi/512
  assign sin[47]  =  8'b11101110;     //47pi/512
  assign cos[47]  =  8'b00111101;     //47pi/512
  assign sin[48]  =  8'b11101101;     //48pi/512
  assign cos[48]  =  8'b00111101;     //48pi/512
  assign sin[49]  =  8'b11101101;     //49pi/512
  assign cos[49]  =  8'b00111101;     //49pi/512
  assign sin[50]  =  8'b11101101;     //50pi/512
  assign cos[50]  =  8'b00111101;     //50pi/512
  assign sin[51]  =  8'b11101100;     //51pi/512
  assign cos[51]  =  8'b00111100;     //51pi/512
  assign sin[52]  =  8'b11101100;     //52pi/512
  assign cos[52]  =  8'b00111100;     //52pi/512
  assign sin[53]  =  8'b11101100;     //53pi/512
  assign cos[53]  =  8'b00111100;     //53pi/512
  assign sin[54]  =  8'b11101011;     //54pi/512
  assign cos[54]  =  8'b00111100;     //54pi/512
  assign sin[55]  =  8'b11101011;     //55pi/512
  assign cos[55]  =  8'b00111100;     //55pi/512
  assign sin[56]  =  8'b11101010;     //56pi/512
  assign cos[56]  =  8'b00111100;     //56pi/512
  assign sin[57]  =  8'b11101010;     //57pi/512
  assign cos[57]  =  8'b00111100;     //57pi/512
  assign sin[58]  =  8'b11101010;     //58pi/512
  assign cos[58]  =  8'b00111011;     //58pi/512
  assign sin[59]  =  8'b11101001;     //59pi/512
  assign cos[59]  =  8'b00111011;     //59pi/512
  assign sin[60]  =  8'b11101001;     //60pi/512
  assign cos[60]  =  8'b00111011;     //60pi/512
  assign sin[61]  =  8'b11101001;     //61pi/512
  assign cos[61]  =  8'b00111011;     //61pi/512
  assign sin[62]  =  8'b11101000;     //62pi/512
  assign cos[62]  =  8'b00111011;     //62pi/512
  assign sin[63]  =  8'b11101000;     //63pi/512
  assign cos[63]  =  8'b00111011;     //63pi/512
  assign sin[64]  =  8'b11101000;     //64pi/512
  assign cos[64]  =  8'b00111011;     //64pi/512
  assign sin[65]  =  8'b11100111;     //65pi/512
  assign cos[65]  =  8'b00111010;     //65pi/512
  assign sin[66]  =  8'b11100111;     //66pi/512
  assign cos[66]  =  8'b00111010;     //66pi/512
  assign sin[67]  =  8'b11100110;     //67pi/512
  assign cos[67]  =  8'b00111010;     //67pi/512
  assign sin[68]  =  8'b11100110;     //68pi/512
  assign cos[68]  =  8'b00111010;     //68pi/512
  assign sin[69]  =  8'b11100110;     //69pi/512
  assign cos[69]  =  8'b00111010;     //69pi/512
  assign sin[70]  =  8'b11100101;     //70pi/512
  assign cos[70]  =  8'b00111010;     //70pi/512
  assign sin[71]  =  8'b11100101;     //71pi/512
  assign cos[71]  =  8'b00111010;     //71pi/512
  assign sin[72]  =  8'b11100101;     //72pi/512
  assign cos[72]  =  8'b00111001;     //72pi/512
  assign sin[73]  =  8'b11100100;     //73pi/512
  assign cos[73]  =  8'b00111001;     //73pi/512
  assign sin[74]  =  8'b11100100;     //74pi/512
  assign cos[74]  =  8'b00111001;     //74pi/512
  assign sin[75]  =  8'b11100100;     //75pi/512
  assign cos[75]  =  8'b00111001;     //75pi/512
  assign sin[76]  =  8'b11100011;     //76pi/512
  assign cos[76]  =  8'b00111001;     //76pi/512
  assign sin[77]  =  8'b11100011;     //77pi/512
  assign cos[77]  =  8'b00111000;     //77pi/512
  assign sin[78]  =  8'b11100011;     //78pi/512
  assign cos[78]  =  8'b00111000;     //78pi/512
  assign sin[79]  =  8'b11100010;     //79pi/512
  assign cos[79]  =  8'b00111000;     //79pi/512
  assign sin[80]  =  8'b11100010;     //80pi/512
  assign cos[80]  =  8'b00111000;     //80pi/512
  assign sin[81]  =  8'b11100001;     //81pi/512
  assign cos[81]  =  8'b00111000;     //81pi/512
  assign sin[82]  =  8'b11100001;     //82pi/512
  assign cos[82]  =  8'b00111000;     //82pi/512
  assign sin[83]  =  8'b11100001;     //83pi/512
  assign cos[83]  =  8'b00110111;     //83pi/512
  assign sin[84]  =  8'b11100000;     //84pi/512
  assign cos[84]  =  8'b00110111;     //84pi/512
  assign sin[85]  =  8'b11100000;     //85pi/512
  assign cos[85]  =  8'b00110111;     //85pi/512
  assign sin[86]  =  8'b11100000;     //86pi/512
  assign cos[86]  =  8'b00110111;     //86pi/512
  assign sin[87]  =  8'b11011111;     //87pi/512
  assign cos[87]  =  8'b00110111;     //87pi/512
  assign sin[88]  =  8'b11011111;     //88pi/512
  assign cos[88]  =  8'b00110110;     //88pi/512
  assign sin[89]  =  8'b11011111;     //89pi/512
  assign cos[89]  =  8'b00110110;     //89pi/512
  assign sin[90]  =  8'b11011110;     //90pi/512
  assign cos[90]  =  8'b00110110;     //90pi/512
  assign sin[91]  =  8'b11011110;     //91pi/512
  assign cos[91]  =  8'b00110110;     //91pi/512
  assign sin[92]  =  8'b11011110;     //92pi/512
  assign cos[92]  =  8'b00110110;     //92pi/512
  assign sin[93]  =  8'b11011101;     //93pi/512
  assign cos[93]  =  8'b00110101;     //93pi/512
  assign sin[94]  =  8'b11011101;     //94pi/512
  assign cos[94]  =  8'b00110101;     //94pi/512
  assign sin[95]  =  8'b11011101;     //95pi/512
  assign cos[95]  =  8'b00110101;     //95pi/512
  assign sin[96]  =  8'b11011100;     //96pi/512
  assign cos[96]  =  8'b00110101;     //96pi/512
  assign sin[97]  =  8'b11011100;     //97pi/512
  assign cos[97]  =  8'b00110100;     //97pi/512
  assign sin[98]  =  8'b11011100;     //98pi/512
  assign cos[98]  =  8'b00110100;     //98pi/512
  assign sin[99]  =  8'b11011011;     //99pi/512
  assign cos[99]  =  8'b00110100;     //99pi/512
  assign sin[100]  =  8'b11011011;     //100pi/512
  assign cos[100]  =  8'b00110100;     //100pi/512
  assign sin[101]  =  8'b11011011;     //101pi/512
  assign cos[101]  =  8'b00110100;     //101pi/512
  assign sin[102]  =  8'b11011011;     //102pi/512
  assign cos[102]  =  8'b00110011;     //102pi/512
  assign sin[103]  =  8'b11011010;     //103pi/512
  assign cos[103]  =  8'b00110011;     //103pi/512
  assign sin[104]  =  8'b11011010;     //104pi/512
  assign cos[104]  =  8'b00110011;     //104pi/512
  assign sin[105]  =  8'b11011010;     //105pi/512
  assign cos[105]  =  8'b00110011;     //105pi/512
  assign sin[106]  =  8'b11011001;     //106pi/512
  assign cos[106]  =  8'b00110010;     //106pi/512
  assign sin[107]  =  8'b11011001;     //107pi/512
  assign cos[107]  =  8'b00110010;     //107pi/512
  assign sin[108]  =  8'b11011001;     //108pi/512
  assign cos[108]  =  8'b00110010;     //108pi/512
  assign sin[109]  =  8'b11011000;     //109pi/512
  assign cos[109]  =  8'b00110010;     //109pi/512
  assign sin[110]  =  8'b11011000;     //110pi/512
  assign cos[110]  =  8'b00110001;     //110pi/512
  assign sin[111]  =  8'b11011000;     //111pi/512
  assign cos[111]  =  8'b00110001;     //111pi/512
  assign sin[112]  =  8'b11010111;     //112pi/512
  assign cos[112]  =  8'b00110001;     //112pi/512
  assign sin[113]  =  8'b11010111;     //113pi/512
  assign cos[113]  =  8'b00110001;     //113pi/512
  assign sin[114]  =  8'b11010111;     //114pi/512
  assign cos[114]  =  8'b00110000;     //114pi/512
  assign sin[115]  =  8'b11010110;     //115pi/512
  assign cos[115]  =  8'b00110000;     //115pi/512
  assign sin[116]  =  8'b11010110;     //116pi/512
  assign cos[116]  =  8'b00110000;     //116pi/512
  assign sin[117]  =  8'b11010110;     //117pi/512
  assign cos[117]  =  8'b00110000;     //117pi/512
  assign sin[118]  =  8'b11010110;     //118pi/512
  assign cos[118]  =  8'b00101111;     //118pi/512
  assign sin[119]  =  8'b11010101;     //119pi/512
  assign cos[119]  =  8'b00101111;     //119pi/512
  assign sin[120]  =  8'b11010101;     //120pi/512
  assign cos[120]  =  8'b00101111;     //120pi/512
  assign sin[121]  =  8'b11010101;     //121pi/512
  assign cos[121]  =  8'b00101111;     //121pi/512
  assign sin[122]  =  8'b11010100;     //122pi/512
  assign cos[122]  =  8'b00101110;     //122pi/512
  assign sin[123]  =  8'b11010100;     //123pi/512
  assign cos[123]  =  8'b00101110;     //123pi/512
  assign sin[124]  =  8'b11010100;     //124pi/512
  assign cos[124]  =  8'b00101110;     //124pi/512
  assign sin[125]  =  8'b11010100;     //125pi/512
  assign cos[125]  =  8'b00101110;     //125pi/512
  assign sin[126]  =  8'b11010011;     //126pi/512
  assign cos[126]  =  8'b00101101;     //126pi/512
  assign sin[127]  =  8'b11010011;     //127pi/512
  assign cos[127]  =  8'b00101101;     //127pi/512
  assign sin[128]  =  8'b11010011;     //128pi/512
  assign cos[128]  =  8'b00101101;     //128pi/512
  assign sin[129]  =  8'b11010010;     //129pi/512
  assign cos[129]  =  8'b00101100;     //129pi/512
  assign sin[130]  =  8'b11010010;     //130pi/512
  assign cos[130]  =  8'b00101100;     //130pi/512
  assign sin[131]  =  8'b11010010;     //131pi/512
  assign cos[131]  =  8'b00101100;     //131pi/512
  assign sin[132]  =  8'b11010010;     //132pi/512
  assign cos[132]  =  8'b00101100;     //132pi/512
  assign sin[133]  =  8'b11010001;     //133pi/512
  assign cos[133]  =  8'b00101011;     //133pi/512
  assign sin[134]  =  8'b11010001;     //134pi/512
  assign cos[134]  =  8'b00101011;     //134pi/512
  assign sin[135]  =  8'b11010001;     //135pi/512
  assign cos[135]  =  8'b00101011;     //135pi/512
  assign sin[136]  =  8'b11010001;     //136pi/512
  assign cos[136]  =  8'b00101010;     //136pi/512
  assign sin[137]  =  8'b11010000;     //137pi/512
  assign cos[137]  =  8'b00101010;     //137pi/512
  assign sin[138]  =  8'b11010000;     //138pi/512
  assign cos[138]  =  8'b00101010;     //138pi/512
  assign sin[139]  =  8'b11010000;     //139pi/512
  assign cos[139]  =  8'b00101010;     //139pi/512
  assign sin[140]  =  8'b11010000;     //140pi/512
  assign cos[140]  =  8'b00101001;     //140pi/512
  assign sin[141]  =  8'b11001111;     //141pi/512
  assign cos[141]  =  8'b00101001;     //141pi/512
  assign sin[142]  =  8'b11001111;     //142pi/512
  assign cos[142]  =  8'b00101001;     //142pi/512
  assign sin[143]  =  8'b11001111;     //143pi/512
  assign cos[143]  =  8'b00101000;     //143pi/512
  assign sin[144]  =  8'b11001111;     //144pi/512
  assign cos[144]  =  8'b00101000;     //144pi/512
  assign sin[145]  =  8'b11001110;     //145pi/512
  assign cos[145]  =  8'b00101000;     //145pi/512
  assign sin[146]  =  8'b11001110;     //146pi/512
  assign cos[146]  =  8'b00100111;     //146pi/512
  assign sin[147]  =  8'b11001110;     //147pi/512
  assign cos[147]  =  8'b00100111;     //147pi/512
  assign sin[148]  =  8'b11001110;     //148pi/512
  assign cos[148]  =  8'b00100111;     //148pi/512
  assign sin[149]  =  8'b11001101;     //149pi/512
  assign cos[149]  =  8'b00100111;     //149pi/512
  assign sin[150]  =  8'b11001101;     //150pi/512
  assign cos[150]  =  8'b00100110;     //150pi/512
  assign sin[151]  =  8'b11001101;     //151pi/512
  assign cos[151]  =  8'b00100110;     //151pi/512
  assign sin[152]  =  8'b11001101;     //152pi/512
  assign cos[152]  =  8'b00100110;     //152pi/512
  assign sin[153]  =  8'b11001100;     //153pi/512
  assign cos[153]  =  8'b00100101;     //153pi/512
  assign sin[154]  =  8'b11001100;     //154pi/512
  assign cos[154]  =  8'b00100101;     //154pi/512
  assign sin[155]  =  8'b11001100;     //155pi/512
  assign cos[155]  =  8'b00100101;     //155pi/512
  assign sin[156]  =  8'b11001100;     //156pi/512
  assign cos[156]  =  8'b00100100;     //156pi/512
  assign sin[157]  =  8'b11001011;     //157pi/512
  assign cos[157]  =  8'b00100100;     //157pi/512
  assign sin[158]  =  8'b11001011;     //158pi/512
  assign cos[158]  =  8'b00100100;     //158pi/512
  assign sin[159]  =  8'b11001011;     //159pi/512
  assign cos[159]  =  8'b00100011;     //159pi/512
  assign sin[160]  =  8'b11001011;     //160pi/512
  assign cos[160]  =  8'b00100011;     //160pi/512
  assign sin[161]  =  8'b11001011;     //161pi/512
  assign cos[161]  =  8'b00100011;     //161pi/512
  assign sin[162]  =  8'b11001010;     //162pi/512
  assign cos[162]  =  8'b00100010;     //162pi/512
  assign sin[163]  =  8'b11001010;     //163pi/512
  assign cos[163]  =  8'b00100010;     //163pi/512
  assign sin[164]  =  8'b11001010;     //164pi/512
  assign cos[164]  =  8'b00100010;     //164pi/512
  assign sin[165]  =  8'b11001010;     //165pi/512
  assign cos[165]  =  8'b00100001;     //165pi/512
  assign sin[166]  =  8'b11001010;     //166pi/512
  assign cos[166]  =  8'b00100001;     //166pi/512
  assign sin[167]  =  8'b11001001;     //167pi/512
  assign cos[167]  =  8'b00100001;     //167pi/512
  assign sin[168]  =  8'b11001001;     //168pi/512
  assign cos[168]  =  8'b00100000;     //168pi/512
  assign sin[169]  =  8'b11001001;     //169pi/512
  assign cos[169]  =  8'b00100000;     //169pi/512
  assign sin[170]  =  8'b11001001;     //170pi/512
  assign cos[170]  =  8'b00100000;     //170pi/512
  assign sin[171]  =  8'b11001001;     //171pi/512
  assign cos[171]  =  8'b00011111;     //171pi/512
  assign sin[172]  =  8'b11001000;     //172pi/512
  assign cos[172]  =  8'b00011111;     //172pi/512
  assign sin[173]  =  8'b11001000;     //173pi/512
  assign cos[173]  =  8'b00011111;     //173pi/512
  assign sin[174]  =  8'b11001000;     //174pi/512
  assign cos[174]  =  8'b00011110;     //174pi/512
  assign sin[175]  =  8'b11001000;     //175pi/512
  assign cos[175]  =  8'b00011110;     //175pi/512
  assign sin[176]  =  8'b11001000;     //176pi/512
  assign cos[176]  =  8'b00011110;     //176pi/512
  assign sin[177]  =  8'b11000111;     //177pi/512
  assign cos[177]  =  8'b00011101;     //177pi/512
  assign sin[178]  =  8'b11000111;     //178pi/512
  assign cos[178]  =  8'b00011101;     //178pi/512
  assign sin[179]  =  8'b11000111;     //179pi/512
  assign cos[179]  =  8'b00011101;     //179pi/512
  assign sin[180]  =  8'b11000111;     //180pi/512
  assign cos[180]  =  8'b00011100;     //180pi/512
  assign sin[181]  =  8'b11000111;     //181pi/512
  assign cos[181]  =  8'b00011100;     //181pi/512
  assign sin[182]  =  8'b11000110;     //182pi/512
  assign cos[182]  =  8'b00011100;     //182pi/512
  assign sin[183]  =  8'b11000110;     //183pi/512
  assign cos[183]  =  8'b00011011;     //183pi/512
  assign sin[184]  =  8'b11000110;     //184pi/512
  assign cos[184]  =  8'b00011011;     //184pi/512
  assign sin[185]  =  8'b11000110;     //185pi/512
  assign cos[185]  =  8'b00011011;     //185pi/512
  assign sin[186]  =  8'b11000110;     //186pi/512
  assign cos[186]  =  8'b00011010;     //186pi/512
  assign sin[187]  =  8'b11000110;     //187pi/512
  assign cos[187]  =  8'b00011010;     //187pi/512
  assign sin[188]  =  8'b11000101;     //188pi/512
  assign cos[188]  =  8'b00011001;     //188pi/512
  assign sin[189]  =  8'b11000101;     //189pi/512
  assign cos[189]  =  8'b00011001;     //189pi/512
  assign sin[190]  =  8'b11000101;     //190pi/512
  assign cos[190]  =  8'b00011001;     //190pi/512
  assign sin[191]  =  8'b11000101;     //191pi/512
  assign cos[191]  =  8'b00011000;     //191pi/512
  assign sin[192]  =  8'b11000101;     //192pi/512
  assign cos[192]  =  8'b00011000;     //192pi/512
  assign sin[193]  =  8'b11000101;     //193pi/512
  assign cos[193]  =  8'b00011000;     //193pi/512
  assign sin[194]  =  8'b11000101;     //194pi/512
  assign cos[194]  =  8'b00010111;     //194pi/512
  assign sin[195]  =  8'b11000100;     //195pi/512
  assign cos[195]  =  8'b00010111;     //195pi/512
  assign sin[196]  =  8'b11000100;     //196pi/512
  assign cos[196]  =  8'b00010111;     //196pi/512
  assign sin[197]  =  8'b11000100;     //197pi/512
  assign cos[197]  =  8'b00010110;     //197pi/512
  assign sin[198]  =  8'b11000100;     //198pi/512
  assign cos[198]  =  8'b00010110;     //198pi/512
  assign sin[199]  =  8'b11000100;     //199pi/512
  assign cos[199]  =  8'b00010101;     //199pi/512
  assign sin[200]  =  8'b11000100;     //200pi/512
  assign cos[200]  =  8'b00010101;     //200pi/512
  assign sin[201]  =  8'b11000100;     //201pi/512
  assign cos[201]  =  8'b00010101;     //201pi/512
  assign sin[202]  =  8'b11000011;     //202pi/512
  assign cos[202]  =  8'b00010100;     //202pi/512
  assign sin[203]  =  8'b11000011;     //203pi/512
  assign cos[203]  =  8'b00010100;     //203pi/512
  assign sin[204]  =  8'b11000011;     //204pi/512
  assign cos[204]  =  8'b00010100;     //204pi/512
  assign sin[205]  =  8'b11000011;     //205pi/512
  assign cos[205]  =  8'b00010011;     //205pi/512
  assign sin[206]  =  8'b11000011;     //206pi/512
  assign cos[206]  =  8'b00010011;     //206pi/512
  assign sin[207]  =  8'b11000011;     //207pi/512
  assign cos[207]  =  8'b00010010;     //207pi/512
  assign sin[208]  =  8'b11000011;     //208pi/512
  assign cos[208]  =  8'b00010010;     //208pi/512
  assign sin[209]  =  8'b11000011;     //209pi/512
  assign cos[209]  =  8'b00010010;     //209pi/512
  assign sin[210]  =  8'b11000011;     //210pi/512
  assign cos[210]  =  8'b00010001;     //210pi/512
  assign sin[211]  =  8'b11000010;     //211pi/512
  assign cos[211]  =  8'b00010001;     //211pi/512
  assign sin[212]  =  8'b11000010;     //212pi/512
  assign cos[212]  =  8'b00010001;     //212pi/512
  assign sin[213]  =  8'b11000010;     //213pi/512
  assign cos[213]  =  8'b00010000;     //213pi/512
  assign sin[214]  =  8'b11000010;     //214pi/512
  assign cos[214]  =  8'b00010000;     //214pi/512
  assign sin[215]  =  8'b11000010;     //215pi/512
  assign cos[215]  =  8'b00001111;     //215pi/512
  assign sin[216]  =  8'b11000010;     //216pi/512
  assign cos[216]  =  8'b00001111;     //216pi/512
  assign sin[217]  =  8'b11000010;     //217pi/512
  assign cos[217]  =  8'b00001111;     //217pi/512
  assign sin[218]  =  8'b11000010;     //218pi/512
  assign cos[218]  =  8'b00001110;     //218pi/512
  assign sin[219]  =  8'b11000010;     //219pi/512
  assign cos[219]  =  8'b00001110;     //219pi/512
  assign sin[220]  =  8'b11000010;     //220pi/512
  assign cos[220]  =  8'b00001110;     //220pi/512
  assign sin[221]  =  8'b11000001;     //221pi/512
  assign cos[221]  =  8'b00001101;     //221pi/512
  assign sin[222]  =  8'b11000001;     //222pi/512
  assign cos[222]  =  8'b00001101;     //222pi/512
  assign sin[223]  =  8'b11000001;     //223pi/512
  assign cos[223]  =  8'b00001100;     //223pi/512
  assign sin[224]  =  8'b11000001;     //224pi/512
  assign cos[224]  =  8'b00001100;     //224pi/512
  assign sin[225]  =  8'b11000001;     //225pi/512
  assign cos[225]  =  8'b00001100;     //225pi/512
  assign sin[226]  =  8'b11000001;     //226pi/512
  assign cos[226]  =  8'b00001011;     //226pi/512
  assign sin[227]  =  8'b11000001;     //227pi/512
  assign cos[227]  =  8'b00001011;     //227pi/512
  assign sin[228]  =  8'b11000001;     //228pi/512
  assign cos[228]  =  8'b00001010;     //228pi/512
  assign sin[229]  =  8'b11000001;     //229pi/512
  assign cos[229]  =  8'b00001010;     //229pi/512
  assign sin[230]  =  8'b11000001;     //230pi/512
  assign cos[230]  =  8'b00001010;     //230pi/512
  assign sin[231]  =  8'b11000001;     //231pi/512
  assign cos[231]  =  8'b00001001;     //231pi/512
  assign sin[232]  =  8'b11000001;     //232pi/512
  assign cos[232]  =  8'b00001001;     //232pi/512
  assign sin[233]  =  8'b11000001;     //233pi/512
  assign cos[233]  =  8'b00001001;     //233pi/512
  assign sin[234]  =  8'b11000001;     //234pi/512
  assign cos[234]  =  8'b00001000;     //234pi/512
  assign sin[235]  =  8'b11000001;     //235pi/512
  assign cos[235]  =  8'b00001000;     //235pi/512
  assign sin[236]  =  8'b11000000;     //236pi/512
  assign cos[236]  =  8'b00000111;     //236pi/512
  assign sin[237]  =  8'b11000000;     //237pi/512
  assign cos[237]  =  8'b00000111;     //237pi/512
  assign sin[238]  =  8'b11000000;     //238pi/512
  assign cos[238]  =  8'b00000111;     //238pi/512
  assign sin[239]  =  8'b11000000;     //239pi/512
  assign cos[239]  =  8'b00000110;     //239pi/512
  assign sin[240]  =  8'b11000000;     //240pi/512
  assign cos[240]  =  8'b00000110;     //240pi/512
  assign sin[241]  =  8'b11000000;     //241pi/512
  assign cos[241]  =  8'b00000101;     //241pi/512
  assign sin[242]  =  8'b11000000;     //242pi/512
  assign cos[242]  =  8'b00000101;     //242pi/512
  assign sin[243]  =  8'b11000000;     //243pi/512
  assign cos[243]  =  8'b00000101;     //243pi/512
  assign sin[244]  =  8'b11000000;     //244pi/512
  assign cos[244]  =  8'b00000100;     //244pi/512
  assign sin[245]  =  8'b11000000;     //245pi/512
  assign cos[245]  =  8'b00000100;     //245pi/512
  assign sin[246]  =  8'b11000000;     //246pi/512
  assign cos[246]  =  8'b00000011;     //246pi/512
  assign sin[247]  =  8'b11000000;     //247pi/512
  assign cos[247]  =  8'b00000011;     //247pi/512
  assign sin[248]  =  8'b11000000;     //248pi/512
  assign cos[248]  =  8'b00000011;     //248pi/512
  assign sin[249]  =  8'b11000000;     //249pi/512
  assign cos[249]  =  8'b00000010;     //249pi/512
  assign sin[250]  =  8'b11000000;     //250pi/512
  assign cos[250]  =  8'b00000010;     //250pi/512
  assign sin[251]  =  8'b11000000;     //251pi/512
  assign cos[251]  =  8'b00000001;     //251pi/512
  assign sin[252]  =  8'b11000000;     //252pi/512
  assign cos[252]  =  8'b00000001;     //252pi/512
  assign sin[253]  =  8'b11000000;     //253pi/512
  assign cos[253]  =  8'b00000001;     //253pi/512
  assign sin[254]  =  8'b11000000;     //254pi/512
  assign cos[254]  =  8'b00000000;     //254pi/512
  assign sin[255]  =  8'b11000000;     //255pi/512
  assign cos[255]  =  8'b00000000;     //255pi/512
  assign sin[256]  =  8'b11000000;     //256pi/512
  assign cos[256]  =  8'b00000000;     //256pi/512
  assign sin[257]  =  8'b11000000;     //257pi/512
  assign cos[257]  =  8'b00000000;     //257pi/512
  assign sin[258]  =  8'b11000000;     //258pi/512
  assign cos[258]  =  8'b11111111;     //258pi/512
  assign sin[259]  =  8'b11000000;     //259pi/512
  assign cos[259]  =  8'b11111111;     //259pi/512
  assign sin[260]  =  8'b11000000;     //260pi/512
  assign cos[260]  =  8'b11111110;     //260pi/512
  assign sin[261]  =  8'b11000000;     //261pi/512
  assign cos[261]  =  8'b11111110;     //261pi/512
  assign sin[262]  =  8'b11000000;     //262pi/512
  assign cos[262]  =  8'b11111110;     //262pi/512
  assign sin[263]  =  8'b11000000;     //263pi/512
  assign cos[263]  =  8'b11111101;     //263pi/512
  assign sin[264]  =  8'b11000000;     //264pi/512
  assign cos[264]  =  8'b11111101;     //264pi/512
  assign sin[265]  =  8'b11000000;     //265pi/512
  assign cos[265]  =  8'b11111100;     //265pi/512
  assign sin[266]  =  8'b11000000;     //266pi/512
  assign cos[266]  =  8'b11111100;     //266pi/512
  assign sin[267]  =  8'b11000000;     //267pi/512
  assign cos[267]  =  8'b11111100;     //267pi/512
  assign sin[268]  =  8'b11000000;     //268pi/512
  assign cos[268]  =  8'b11111011;     //268pi/512
  assign sin[269]  =  8'b11000000;     //269pi/512
  assign cos[269]  =  8'b11111011;     //269pi/512
  assign sin[270]  =  8'b11000000;     //270pi/512
  assign cos[270]  =  8'b11111011;     //270pi/512
  assign sin[271]  =  8'b11000000;     //271pi/512
  assign cos[271]  =  8'b11111010;     //271pi/512
  assign sin[272]  =  8'b11000000;     //272pi/512
  assign cos[272]  =  8'b11111010;     //272pi/512
  assign sin[273]  =  8'b11000000;     //273pi/512
  assign cos[273]  =  8'b11111001;     //273pi/512
  assign sin[274]  =  8'b11000000;     //274pi/512
  assign cos[274]  =  8'b11111001;     //274pi/512
  assign sin[275]  =  8'b11000000;     //275pi/512
  assign cos[275]  =  8'b11111001;     //275pi/512
  assign sin[276]  =  8'b11000000;     //276pi/512
  assign cos[276]  =  8'b11111000;     //276pi/512
  assign sin[277]  =  8'b11000001;     //277pi/512
  assign cos[277]  =  8'b11111000;     //277pi/512
  assign sin[278]  =  8'b11000001;     //278pi/512
  assign cos[278]  =  8'b11110111;     //278pi/512
  assign sin[279]  =  8'b11000001;     //279pi/512
  assign cos[279]  =  8'b11110111;     //279pi/512
  assign sin[280]  =  8'b11000001;     //280pi/512
  assign cos[280]  =  8'b11110111;     //280pi/512
  assign sin[281]  =  8'b11000001;     //281pi/512
  assign cos[281]  =  8'b11110110;     //281pi/512
  assign sin[282]  =  8'b11000001;     //282pi/512
  assign cos[282]  =  8'b11110110;     //282pi/512
  assign sin[283]  =  8'b11000001;     //283pi/512
  assign cos[283]  =  8'b11110101;     //283pi/512
  assign sin[284]  =  8'b11000001;     //284pi/512
  assign cos[284]  =  8'b11110101;     //284pi/512
  assign sin[285]  =  8'b11000001;     //285pi/512
  assign cos[285]  =  8'b11110101;     //285pi/512
  assign sin[286]  =  8'b11000001;     //286pi/512
  assign cos[286]  =  8'b11110100;     //286pi/512
  assign sin[287]  =  8'b11000001;     //287pi/512
  assign cos[287]  =  8'b11110100;     //287pi/512
  assign sin[288]  =  8'b11000001;     //288pi/512
  assign cos[288]  =  8'b11110100;     //288pi/512
  assign sin[289]  =  8'b11000001;     //289pi/512
  assign cos[289]  =  8'b11110011;     //289pi/512
  assign sin[290]  =  8'b11000001;     //290pi/512
  assign cos[290]  =  8'b11110011;     //290pi/512
  assign sin[291]  =  8'b11000001;     //291pi/512
  assign cos[291]  =  8'b11110010;     //291pi/512
  assign sin[292]  =  8'b11000010;     //292pi/512
  assign cos[292]  =  8'b11110010;     //292pi/512
  assign sin[293]  =  8'b11000010;     //293pi/512
  assign cos[293]  =  8'b11110010;     //293pi/512
  assign sin[294]  =  8'b11000010;     //294pi/512
  assign cos[294]  =  8'b11110001;     //294pi/512
  assign sin[295]  =  8'b11000010;     //295pi/512
  assign cos[295]  =  8'b11110001;     //295pi/512
  assign sin[296]  =  8'b11000010;     //296pi/512
  assign cos[296]  =  8'b11110000;     //296pi/512
  assign sin[297]  =  8'b11000010;     //297pi/512
  assign cos[297]  =  8'b11110000;     //297pi/512
  assign sin[298]  =  8'b11000010;     //298pi/512
  assign cos[298]  =  8'b11110000;     //298pi/512
  assign sin[299]  =  8'b11000010;     //299pi/512
  assign cos[299]  =  8'b11101111;     //299pi/512
  assign sin[300]  =  8'b11000010;     //300pi/512
  assign cos[300]  =  8'b11101111;     //300pi/512
  assign sin[301]  =  8'b11000010;     //301pi/512
  assign cos[301]  =  8'b11101111;     //301pi/512
  assign sin[302]  =  8'b11000011;     //302pi/512
  assign cos[302]  =  8'b11101110;     //302pi/512
  assign sin[303]  =  8'b11000011;     //303pi/512
  assign cos[303]  =  8'b11101110;     //303pi/512
  assign sin[304]  =  8'b11000011;     //304pi/512
  assign cos[304]  =  8'b11101101;     //304pi/512
  assign sin[305]  =  8'b11000011;     //305pi/512
  assign cos[305]  =  8'b11101101;     //305pi/512
  assign sin[306]  =  8'b11000011;     //306pi/512
  assign cos[306]  =  8'b11101101;     //306pi/512
  assign sin[307]  =  8'b11000011;     //307pi/512
  assign cos[307]  =  8'b11101100;     //307pi/512
  assign sin[308]  =  8'b11000011;     //308pi/512
  assign cos[308]  =  8'b11101100;     //308pi/512
  assign sin[309]  =  8'b11000011;     //309pi/512
  assign cos[309]  =  8'b11101100;     //309pi/512
  assign sin[310]  =  8'b11000011;     //310pi/512
  assign cos[310]  =  8'b11101011;     //310pi/512
  assign sin[311]  =  8'b11000100;     //311pi/512
  assign cos[311]  =  8'b11101011;     //311pi/512
  assign sin[312]  =  8'b11000100;     //312pi/512
  assign cos[312]  =  8'b11101010;     //312pi/512
  assign sin[313]  =  8'b11000100;     //313pi/512
  assign cos[313]  =  8'b11101010;     //313pi/512
  assign sin[314]  =  8'b11000100;     //314pi/512
  assign cos[314]  =  8'b11101010;     //314pi/512
  assign sin[315]  =  8'b11000100;     //315pi/512
  assign cos[315]  =  8'b11101001;     //315pi/512
  assign sin[316]  =  8'b11000100;     //316pi/512
  assign cos[316]  =  8'b11101001;     //316pi/512
  assign sin[317]  =  8'b11000100;     //317pi/512
  assign cos[317]  =  8'b11101001;     //317pi/512
  assign sin[318]  =  8'b11000101;     //318pi/512
  assign cos[318]  =  8'b11101000;     //318pi/512
  assign sin[319]  =  8'b11000101;     //319pi/512
  assign cos[319]  =  8'b11101000;     //319pi/512
  assign sin[320]  =  8'b11000101;     //320pi/512
  assign cos[320]  =  8'b11101000;     //320pi/512
  assign sin[321]  =  8'b11000101;     //321pi/512
  assign cos[321]  =  8'b11100111;     //321pi/512
  assign sin[322]  =  8'b11000101;     //322pi/512
  assign cos[322]  =  8'b11100111;     //322pi/512
  assign sin[323]  =  8'b11000101;     //323pi/512
  assign cos[323]  =  8'b11100110;     //323pi/512
  assign sin[324]  =  8'b11000101;     //324pi/512
  assign cos[324]  =  8'b11100110;     //324pi/512
  assign sin[325]  =  8'b11000110;     //325pi/512
  assign cos[325]  =  8'b11100110;     //325pi/512
  assign sin[326]  =  8'b11000110;     //326pi/512
  assign cos[326]  =  8'b11100101;     //326pi/512
  assign sin[327]  =  8'b11000110;     //327pi/512
  assign cos[327]  =  8'b11100101;     //327pi/512
  assign sin[328]  =  8'b11000110;     //328pi/512
  assign cos[328]  =  8'b11100101;     //328pi/512
  assign sin[329]  =  8'b11000110;     //329pi/512
  assign cos[329]  =  8'b11100100;     //329pi/512
  assign sin[330]  =  8'b11000110;     //330pi/512
  assign cos[330]  =  8'b11100100;     //330pi/512
  assign sin[331]  =  8'b11000111;     //331pi/512
  assign cos[331]  =  8'b11100100;     //331pi/512
  assign sin[332]  =  8'b11000111;     //332pi/512
  assign cos[332]  =  8'b11100011;     //332pi/512
  assign sin[333]  =  8'b11000111;     //333pi/512
  assign cos[333]  =  8'b11100011;     //333pi/512
  assign sin[334]  =  8'b11000111;     //334pi/512
  assign cos[334]  =  8'b11100011;     //334pi/512
  assign sin[335]  =  8'b11000111;     //335pi/512
  assign cos[335]  =  8'b11100010;     //335pi/512
  assign sin[336]  =  8'b11001000;     //336pi/512
  assign cos[336]  =  8'b11100010;     //336pi/512
  assign sin[337]  =  8'b11001000;     //337pi/512
  assign cos[337]  =  8'b11100001;     //337pi/512
  assign sin[338]  =  8'b11001000;     //338pi/512
  assign cos[338]  =  8'b11100001;     //338pi/512
  assign sin[339]  =  8'b11001000;     //339pi/512
  assign cos[339]  =  8'b11100001;     //339pi/512
  assign sin[340]  =  8'b11001000;     //340pi/512
  assign cos[340]  =  8'b11100000;     //340pi/512
  assign sin[341]  =  8'b11001001;     //341pi/512
  assign cos[341]  =  8'b11100000;     //341pi/512
  assign sin[342]  =  8'b11001001;     //342pi/512
  assign cos[342]  =  8'b11100000;     //342pi/512
  assign sin[343]  =  8'b11001001;     //343pi/512
  assign cos[343]  =  8'b11011111;     //343pi/512
  assign sin[344]  =  8'b11001001;     //344pi/512
  assign cos[344]  =  8'b11011111;     //344pi/512
  assign sin[345]  =  8'b11001001;     //345pi/512
  assign cos[345]  =  8'b11011111;     //345pi/512
  assign sin[346]  =  8'b11001010;     //346pi/512
  assign cos[346]  =  8'b11011110;     //346pi/512
  assign sin[347]  =  8'b11001010;     //347pi/512
  assign cos[347]  =  8'b11011110;     //347pi/512
  assign sin[348]  =  8'b11001010;     //348pi/512
  assign cos[348]  =  8'b11011110;     //348pi/512
  assign sin[349]  =  8'b11001010;     //349pi/512
  assign cos[349]  =  8'b11011101;     //349pi/512
  assign sin[350]  =  8'b11001010;     //350pi/512
  assign cos[350]  =  8'b11011101;     //350pi/512
  assign sin[351]  =  8'b11001011;     //351pi/512
  assign cos[351]  =  8'b11011101;     //351pi/512
  assign sin[352]  =  8'b11001011;     //352pi/512
  assign cos[352]  =  8'b11011100;     //352pi/512
  assign sin[353]  =  8'b11001011;     //353pi/512
  assign cos[353]  =  8'b11011100;     //353pi/512
  assign sin[354]  =  8'b11001011;     //354pi/512
  assign cos[354]  =  8'b11011100;     //354pi/512
  assign sin[355]  =  8'b11001011;     //355pi/512
  assign cos[355]  =  8'b11011011;     //355pi/512
  assign sin[356]  =  8'b11001100;     //356pi/512
  assign cos[356]  =  8'b11011011;     //356pi/512
  assign sin[357]  =  8'b11001100;     //357pi/512
  assign cos[357]  =  8'b11011011;     //357pi/512
  assign sin[358]  =  8'b11001100;     //358pi/512
  assign cos[358]  =  8'b11011011;     //358pi/512
  assign sin[359]  =  8'b11001100;     //359pi/512
  assign cos[359]  =  8'b11011010;     //359pi/512
  assign sin[360]  =  8'b11001101;     //360pi/512
  assign cos[360]  =  8'b11011010;     //360pi/512
  assign sin[361]  =  8'b11001101;     //361pi/512
  assign cos[361]  =  8'b11011010;     //361pi/512
  assign sin[362]  =  8'b11001101;     //362pi/512
  assign cos[362]  =  8'b11011001;     //362pi/512
  assign sin[363]  =  8'b11001101;     //363pi/512
  assign cos[363]  =  8'b11011001;     //363pi/512
  assign sin[364]  =  8'b11001110;     //364pi/512
  assign cos[364]  =  8'b11011001;     //364pi/512
  assign sin[365]  =  8'b11001110;     //365pi/512
  assign cos[365]  =  8'b11011000;     //365pi/512
  assign sin[366]  =  8'b11001110;     //366pi/512
  assign cos[366]  =  8'b11011000;     //366pi/512
  assign sin[367]  =  8'b11001110;     //367pi/512
  assign cos[367]  =  8'b11011000;     //367pi/512
  assign sin[368]  =  8'b11001111;     //368pi/512
  assign cos[368]  =  8'b11010111;     //368pi/512
  assign sin[369]  =  8'b11001111;     //369pi/512
  assign cos[369]  =  8'b11010111;     //369pi/512
  assign sin[370]  =  8'b11001111;     //370pi/512
  assign cos[370]  =  8'b11010111;     //370pi/512
  assign sin[371]  =  8'b11001111;     //371pi/512
  assign cos[371]  =  8'b11010110;     //371pi/512
  assign sin[372]  =  8'b11010000;     //372pi/512
  assign cos[372]  =  8'b11010110;     //372pi/512
  assign sin[373]  =  8'b11010000;     //373pi/512
  assign cos[373]  =  8'b11010110;     //373pi/512
  assign sin[374]  =  8'b11010000;     //374pi/512
  assign cos[374]  =  8'b11010110;     //374pi/512
  assign sin[375]  =  8'b11010000;     //375pi/512
  assign cos[375]  =  8'b11010101;     //375pi/512
  assign sin[376]  =  8'b11010001;     //376pi/512
  assign cos[376]  =  8'b11010101;     //376pi/512
  assign sin[377]  =  8'b11010001;     //377pi/512
  assign cos[377]  =  8'b11010101;     //377pi/512
  assign sin[378]  =  8'b11010001;     //378pi/512
  assign cos[378]  =  8'b11010100;     //378pi/512
  assign sin[379]  =  8'b11010001;     //379pi/512
  assign cos[379]  =  8'b11010100;     //379pi/512
  assign sin[380]  =  8'b11010010;     //380pi/512
  assign cos[380]  =  8'b11010100;     //380pi/512
  assign sin[381]  =  8'b11010010;     //381pi/512
  assign cos[381]  =  8'b11010100;     //381pi/512
  assign sin[382]  =  8'b11010010;     //382pi/512
  assign cos[382]  =  8'b11010011;     //382pi/512
  assign sin[383]  =  8'b11010010;     //383pi/512
  assign cos[383]  =  8'b11010011;     //383pi/512
  assign sin[384]  =  8'b11010011;     //384pi/512
  assign cos[384]  =  8'b11010011;     //384pi/512
  assign sin[385]  =  8'b11010011;     //385pi/512
  assign cos[385]  =  8'b11010010;     //385pi/512
  assign sin[386]  =  8'b11010011;     //386pi/512
  assign cos[386]  =  8'b11010010;     //386pi/512
  assign sin[387]  =  8'b11010100;     //387pi/512
  assign cos[387]  =  8'b11010010;     //387pi/512
  assign sin[388]  =  8'b11010100;     //388pi/512
  assign cos[388]  =  8'b11010010;     //388pi/512
  assign sin[389]  =  8'b11010100;     //389pi/512
  assign cos[389]  =  8'b11010001;     //389pi/512
  assign sin[390]  =  8'b11010100;     //390pi/512
  assign cos[390]  =  8'b11010001;     //390pi/512
  assign sin[391]  =  8'b11010101;     //391pi/512
  assign cos[391]  =  8'b11010001;     //391pi/512
  assign sin[392]  =  8'b11010101;     //392pi/512
  assign cos[392]  =  8'b11010001;     //392pi/512
  assign sin[393]  =  8'b11010101;     //393pi/512
  assign cos[393]  =  8'b11010000;     //393pi/512
  assign sin[394]  =  8'b11010110;     //394pi/512
  assign cos[394]  =  8'b11010000;     //394pi/512
  assign sin[395]  =  8'b11010110;     //395pi/512
  assign cos[395]  =  8'b11010000;     //395pi/512
  assign sin[396]  =  8'b11010110;     //396pi/512
  assign cos[396]  =  8'b11010000;     //396pi/512
  assign sin[397]  =  8'b11010110;     //397pi/512
  assign cos[397]  =  8'b11001111;     //397pi/512
  assign sin[398]  =  8'b11010111;     //398pi/512
  assign cos[398]  =  8'b11001111;     //398pi/512
  assign sin[399]  =  8'b11010111;     //399pi/512
  assign cos[399]  =  8'b11001111;     //399pi/512
  assign sin[400]  =  8'b11010111;     //400pi/512
  assign cos[400]  =  8'b11001111;     //400pi/512
  assign sin[401]  =  8'b11011000;     //401pi/512
  assign cos[401]  =  8'b11001110;     //401pi/512
  assign sin[402]  =  8'b11011000;     //402pi/512
  assign cos[402]  =  8'b11001110;     //402pi/512
  assign sin[403]  =  8'b11011000;     //403pi/512
  assign cos[403]  =  8'b11001110;     //403pi/512
  assign sin[404]  =  8'b11011001;     //404pi/512
  assign cos[404]  =  8'b11001110;     //404pi/512
  assign sin[405]  =  8'b11011001;     //405pi/512
  assign cos[405]  =  8'b11001101;     //405pi/512
  assign sin[406]  =  8'b11011001;     //406pi/512
  assign cos[406]  =  8'b11001101;     //406pi/512
  assign sin[407]  =  8'b11011010;     //407pi/512
  assign cos[407]  =  8'b11001101;     //407pi/512
  assign sin[408]  =  8'b11011010;     //408pi/512
  assign cos[408]  =  8'b11001101;     //408pi/512
  assign sin[409]  =  8'b11011010;     //409pi/512
  assign cos[409]  =  8'b11001100;     //409pi/512
  assign sin[410]  =  8'b11011011;     //410pi/512
  assign cos[410]  =  8'b11001100;     //410pi/512
  assign sin[411]  =  8'b11011011;     //411pi/512
  assign cos[411]  =  8'b11001100;     //411pi/512
  assign sin[412]  =  8'b11011011;     //412pi/512
  assign cos[412]  =  8'b11001100;     //412pi/512
  assign sin[413]  =  8'b11011011;     //413pi/512
  assign cos[413]  =  8'b11001011;     //413pi/512
  assign sin[414]  =  8'b11011100;     //414pi/512
  assign cos[414]  =  8'b11001011;     //414pi/512
  assign sin[415]  =  8'b11011100;     //415pi/512
  assign cos[415]  =  8'b11001011;     //415pi/512
  assign sin[416]  =  8'b11011100;     //416pi/512
  assign cos[416]  =  8'b11001011;     //416pi/512
  assign sin[417]  =  8'b11011101;     //417pi/512
  assign cos[417]  =  8'b11001011;     //417pi/512
  assign sin[418]  =  8'b11011101;     //418pi/512
  assign cos[418]  =  8'b11001010;     //418pi/512
  assign sin[419]  =  8'b11011101;     //419pi/512
  assign cos[419]  =  8'b11001010;     //419pi/512
  assign sin[420]  =  8'b11011110;     //420pi/512
  assign cos[420]  =  8'b11001010;     //420pi/512
  assign sin[421]  =  8'b11011110;     //421pi/512
  assign cos[421]  =  8'b11001010;     //421pi/512
  assign sin[422]  =  8'b11011110;     //422pi/512
  assign cos[422]  =  8'b11001010;     //422pi/512
  assign sin[423]  =  8'b11011111;     //423pi/512
  assign cos[423]  =  8'b11001001;     //423pi/512
  assign sin[424]  =  8'b11011111;     //424pi/512
  assign cos[424]  =  8'b11001001;     //424pi/512
  assign sin[425]  =  8'b11011111;     //425pi/512
  assign cos[425]  =  8'b11001001;     //425pi/512
  assign sin[426]  =  8'b11100000;     //426pi/512
  assign cos[426]  =  8'b11001001;     //426pi/512
  assign sin[427]  =  8'b11100000;     //427pi/512
  assign cos[427]  =  8'b11001001;     //427pi/512
  assign sin[428]  =  8'b11100000;     //428pi/512
  assign cos[428]  =  8'b11001000;     //428pi/512
  assign sin[429]  =  8'b11100001;     //429pi/512
  assign cos[429]  =  8'b11001000;     //429pi/512
  assign sin[430]  =  8'b11100001;     //430pi/512
  assign cos[430]  =  8'b11001000;     //430pi/512
  assign sin[431]  =  8'b11100001;     //431pi/512
  assign cos[431]  =  8'b11001000;     //431pi/512
  assign sin[432]  =  8'b11100010;     //432pi/512
  assign cos[432]  =  8'b11001000;     //432pi/512
  assign sin[433]  =  8'b11100010;     //433pi/512
  assign cos[433]  =  8'b11000111;     //433pi/512
  assign sin[434]  =  8'b11100011;     //434pi/512
  assign cos[434]  =  8'b11000111;     //434pi/512
  assign sin[435]  =  8'b11100011;     //435pi/512
  assign cos[435]  =  8'b11000111;     //435pi/512
  assign sin[436]  =  8'b11100011;     //436pi/512
  assign cos[436]  =  8'b11000111;     //436pi/512
  assign sin[437]  =  8'b11100100;     //437pi/512
  assign cos[437]  =  8'b11000111;     //437pi/512
  assign sin[438]  =  8'b11100100;     //438pi/512
  assign cos[438]  =  8'b11000110;     //438pi/512
  assign sin[439]  =  8'b11100100;     //439pi/512
  assign cos[439]  =  8'b11000110;     //439pi/512
  assign sin[440]  =  8'b11100101;     //440pi/512
  assign cos[440]  =  8'b11000110;     //440pi/512
  assign sin[441]  =  8'b11100101;     //441pi/512
  assign cos[441]  =  8'b11000110;     //441pi/512
  assign sin[442]  =  8'b11100101;     //442pi/512
  assign cos[442]  =  8'b11000110;     //442pi/512
  assign sin[443]  =  8'b11100110;     //443pi/512
  assign cos[443]  =  8'b11000110;     //443pi/512
  assign sin[444]  =  8'b11100110;     //444pi/512
  assign cos[444]  =  8'b11000101;     //444pi/512
  assign sin[445]  =  8'b11100110;     //445pi/512
  assign cos[445]  =  8'b11000101;     //445pi/512
  assign sin[446]  =  8'b11100111;     //446pi/512
  assign cos[446]  =  8'b11000101;     //446pi/512
  assign sin[447]  =  8'b11100111;     //447pi/512
  assign cos[447]  =  8'b11000101;     //447pi/512
  assign sin[448]  =  8'b11101000;     //448pi/512
  assign cos[448]  =  8'b11000101;     //448pi/512
  assign sin[449]  =  8'b11101000;     //449pi/512
  assign cos[449]  =  8'b11000101;     //449pi/512
  assign sin[450]  =  8'b11101000;     //450pi/512
  assign cos[450]  =  8'b11000101;     //450pi/512
  assign sin[451]  =  8'b11101001;     //451pi/512
  assign cos[451]  =  8'b11000100;     //451pi/512
  assign sin[452]  =  8'b11101001;     //452pi/512
  assign cos[452]  =  8'b11000100;     //452pi/512
  assign sin[453]  =  8'b11101001;     //453pi/512
  assign cos[453]  =  8'b11000100;     //453pi/512
  assign sin[454]  =  8'b11101010;     //454pi/512
  assign cos[454]  =  8'b11000100;     //454pi/512
  assign sin[455]  =  8'b11101010;     //455pi/512
  assign cos[455]  =  8'b11000100;     //455pi/512
  assign sin[456]  =  8'b11101010;     //456pi/512
  assign cos[456]  =  8'b11000100;     //456pi/512
  assign sin[457]  =  8'b11101011;     //457pi/512
  assign cos[457]  =  8'b11000100;     //457pi/512
  assign sin[458]  =  8'b11101011;     //458pi/512
  assign cos[458]  =  8'b11000011;     //458pi/512
  assign sin[459]  =  8'b11101100;     //459pi/512
  assign cos[459]  =  8'b11000011;     //459pi/512
  assign sin[460]  =  8'b11101100;     //460pi/512
  assign cos[460]  =  8'b11000011;     //460pi/512
  assign sin[461]  =  8'b11101100;     //461pi/512
  assign cos[461]  =  8'b11000011;     //461pi/512
  assign sin[462]  =  8'b11101101;     //462pi/512
  assign cos[462]  =  8'b11000011;     //462pi/512
  assign sin[463]  =  8'b11101101;     //463pi/512
  assign cos[463]  =  8'b11000011;     //463pi/512
  assign sin[464]  =  8'b11101101;     //464pi/512
  assign cos[464]  =  8'b11000011;     //464pi/512
  assign sin[465]  =  8'b11101110;     //465pi/512
  assign cos[465]  =  8'b11000011;     //465pi/512
  assign sin[466]  =  8'b11101110;     //466pi/512
  assign cos[466]  =  8'b11000011;     //466pi/512
  assign sin[467]  =  8'b11101111;     //467pi/512
  assign cos[467]  =  8'b11000010;     //467pi/512
  assign sin[468]  =  8'b11101111;     //468pi/512
  assign cos[468]  =  8'b11000010;     //468pi/512
  assign sin[469]  =  8'b11101111;     //469pi/512
  assign cos[469]  =  8'b11000010;     //469pi/512
  assign sin[470]  =  8'b11110000;     //470pi/512
  assign cos[470]  =  8'b11000010;     //470pi/512
  assign sin[471]  =  8'b11110000;     //471pi/512
  assign cos[471]  =  8'b11000010;     //471pi/512
  assign sin[472]  =  8'b11110000;     //472pi/512
  assign cos[472]  =  8'b11000010;     //472pi/512
  assign sin[473]  =  8'b11110001;     //473pi/512
  assign cos[473]  =  8'b11000010;     //473pi/512
  assign sin[474]  =  8'b11110001;     //474pi/512
  assign cos[474]  =  8'b11000010;     //474pi/512
  assign sin[475]  =  8'b11110010;     //475pi/512
  assign cos[475]  =  8'b11000010;     //475pi/512
  assign sin[476]  =  8'b11110010;     //476pi/512
  assign cos[476]  =  8'b11000010;     //476pi/512
  assign sin[477]  =  8'b11110010;     //477pi/512
  assign cos[477]  =  8'b11000001;     //477pi/512
  assign sin[478]  =  8'b11110011;     //478pi/512
  assign cos[478]  =  8'b11000001;     //478pi/512
  assign sin[479]  =  8'b11110011;     //479pi/512
  assign cos[479]  =  8'b11000001;     //479pi/512
  assign sin[480]  =  8'b11110100;     //480pi/512
  assign cos[480]  =  8'b11000001;     //480pi/512
  assign sin[481]  =  8'b11110100;     //481pi/512
  assign cos[481]  =  8'b11000001;     //481pi/512
  assign sin[482]  =  8'b11110100;     //482pi/512
  assign cos[482]  =  8'b11000001;     //482pi/512
  assign sin[483]  =  8'b11110101;     //483pi/512
  assign cos[483]  =  8'b11000001;     //483pi/512
  assign sin[484]  =  8'b11110101;     //484pi/512
  assign cos[484]  =  8'b11000001;     //484pi/512
  assign sin[485]  =  8'b11110101;     //485pi/512
  assign cos[485]  =  8'b11000001;     //485pi/512
  assign sin[486]  =  8'b11110110;     //486pi/512
  assign cos[486]  =  8'b11000001;     //486pi/512
  assign sin[487]  =  8'b11110110;     //487pi/512
  assign cos[487]  =  8'b11000001;     //487pi/512
  assign sin[488]  =  8'b11110111;     //488pi/512
  assign cos[488]  =  8'b11000001;     //488pi/512
  assign sin[489]  =  8'b11110111;     //489pi/512
  assign cos[489]  =  8'b11000001;     //489pi/512
  assign sin[490]  =  8'b11110111;     //490pi/512
  assign cos[490]  =  8'b11000001;     //490pi/512
  assign sin[491]  =  8'b11111000;     //491pi/512
  assign cos[491]  =  8'b11000001;     //491pi/512
  assign sin[492]  =  8'b11111000;     //492pi/512
  assign cos[492]  =  8'b11000000;     //492pi/512
  assign sin[493]  =  8'b11111001;     //493pi/512
  assign cos[493]  =  8'b11000000;     //493pi/512
  assign sin[494]  =  8'b11111001;     //494pi/512
  assign cos[494]  =  8'b11000000;     //494pi/512
  assign sin[495]  =  8'b11111001;     //495pi/512
  assign cos[495]  =  8'b11000000;     //495pi/512
  assign sin[496]  =  8'b11111010;     //496pi/512
  assign cos[496]  =  8'b11000000;     //496pi/512
  assign sin[497]  =  8'b11111010;     //497pi/512
  assign cos[497]  =  8'b11000000;     //497pi/512
  assign sin[498]  =  8'b11111011;     //498pi/512
  assign cos[498]  =  8'b11000000;     //498pi/512
  assign sin[499]  =  8'b11111011;     //499pi/512
  assign cos[499]  =  8'b11000000;     //499pi/512
  assign sin[500]  =  8'b11111011;     //500pi/512
  assign cos[500]  =  8'b11000000;     //500pi/512
  assign sin[501]  =  8'b11111100;     //501pi/512
  assign cos[501]  =  8'b11000000;     //501pi/512
  assign sin[502]  =  8'b11111100;     //502pi/512
  assign cos[502]  =  8'b11000000;     //502pi/512
  assign sin[503]  =  8'b11111100;     //503pi/512
  assign cos[503]  =  8'b11000000;     //503pi/512
  assign sin[504]  =  8'b11111101;     //504pi/512
  assign cos[504]  =  8'b11000000;     //504pi/512
  assign sin[505]  =  8'b11111101;     //505pi/512
  assign cos[505]  =  8'b11000000;     //505pi/512
  assign sin[506]  =  8'b11111110;     //506pi/512
  assign cos[506]  =  8'b11000000;     //506pi/512
  assign sin[507]  =  8'b11111110;     //507pi/512
  assign cos[507]  =  8'b11000000;     //507pi/512
  assign sin[508]  =  8'b11111110;     //508pi/512
  assign cos[508]  =  8'b11000000;     //508pi/512
  assign sin[509]  =  8'b11111111;     //509pi/512
  assign cos[509]  =  8'b11000000;     //509pi/512
  assign sin[510]  =  8'b11111111;     //510pi/512
  assign cos[510]  =  8'b11000000;     //510pi/512
  assign sin[511]  =  8'b00000000;     //511pi/512
  assign cos[511]  =  8'b11000000;     //511pi/512

endmodule