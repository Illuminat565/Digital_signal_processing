module  M_TWIDLE_15_B_0_20_v  #(parameter SIZE = 10, word_length_tw = 15) (
    input            clk,
    input            en_rd,
    input   [10:0]   rd_ptr_angle,
    input            en_modf,
    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );
reg signed [word_length_tw-1:0]  cos    [511:0];
reg signed [word_length_tw-1:0]  sin    [511:0];
reg signed [word_length_tw-1:0]  m_cos  [511:0];
reg signed [word_length_tw-1:0]  m_sin  [511:0];
reg signed [word_length_tw-1:0]  cos_temp;
reg signed [word_length_tw-1:0]  sin_temp;
reg signed [word_length_tw-1:0]  m_cos_temp;
reg signed [word_length_tw-1:0]  m_sin_temp;
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & ~ en_modf) begin
                  cos_temp           <= cos   [rd_ptr_angle];
                  sin_temp           <= sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & en_modf) begin
                  m_cos_temp           <= m_cos   [rd_ptr_angle];
                  m_sin_temp           <= m_sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(*) begin 
             if (en_modf) begin
                  cos_data           <= m_cos_temp;
                  sin_data           <= m_sin_temp;
             end else begin
                  cos_data           <= cos_temp;
                  sin_data           <= sin_temp;
             end 
        end
initial begin
   sin[0]  =  15'b000000000000000;     //0pi/512
   cos[0]  =  15'b010000000000000;     //0pi/512
   sin[1]  =  15'b111111111001110;     //1pi/512
   cos[1]  =  15'b001111111111111;     //1pi/512
   sin[2]  =  15'b111111110011011;     //2pi/512
   cos[2]  =  15'b001111111111111;     //2pi/512
   sin[3]  =  15'b111111101101001;     //3pi/512
   cos[3]  =  15'b001111111111110;     //3pi/512
   sin[4]  =  15'b111111100110111;     //4pi/512
   cos[4]  =  15'b001111111111101;     //4pi/512
   sin[5]  =  15'b111111100000101;     //5pi/512
   cos[5]  =  15'b001111111111100;     //5pi/512
   sin[6]  =  15'b111111011010010;     //6pi/512
   cos[6]  =  15'b001111111111010;     //6pi/512
   sin[7]  =  15'b111111010100000;     //7pi/512
   cos[7]  =  15'b001111111111000;     //7pi/512
   sin[8]  =  15'b111111001101110;     //8pi/512
   cos[8]  =  15'b001111111110110;     //8pi/512
   sin[9]  =  15'b111111000111100;     //9pi/512
   cos[9]  =  15'b001111111110011;     //9pi/512
   sin[10]  =  15'b111111000001010;     //10pi/512
   cos[10]  =  15'b001111111110000;     //10pi/512
   sin[11]  =  15'b111110111010111;     //11pi/512
   cos[11]  =  15'b001111111101101;     //11pi/512
   sin[12]  =  15'b111110110100101;     //12pi/512
   cos[12]  =  15'b001111111101001;     //12pi/512
   sin[13]  =  15'b111110101110011;     //13pi/512
   cos[13]  =  15'b001111111100101;     //13pi/512
   sin[14]  =  15'b111110101000001;     //14pi/512
   cos[14]  =  15'b001111111100001;     //14pi/512
   sin[15]  =  15'b111110100001111;     //15pi/512
   cos[15]  =  15'b001111111011101;     //15pi/512
   sin[16]  =  15'b111110011011101;     //16pi/512
   cos[16]  =  15'b001111111011000;     //16pi/512
   sin[17]  =  15'b111110010101011;     //17pi/512
   cos[17]  =  15'b001111111010011;     //17pi/512
   sin[18]  =  15'b111110001111001;     //18pi/512
   cos[18]  =  15'b001111111001110;     //18pi/512
   sin[19]  =  15'b111110001000111;     //19pi/512
   cos[19]  =  15'b001111111001000;     //19pi/512
   sin[20]  =  15'b111110000010101;     //20pi/512
   cos[20]  =  15'b001111111000010;     //20pi/512
   sin[21]  =  15'b111101111100011;     //21pi/512
   cos[21]  =  15'b001111110111100;     //21pi/512
   sin[22]  =  15'b111101110110010;     //22pi/512
   cos[22]  =  15'b001111110110101;     //22pi/512
   sin[23]  =  15'b111101110000000;     //23pi/512
   cos[23]  =  15'b001111110101110;     //23pi/512
   sin[24]  =  15'b111101101001110;     //24pi/512
   cos[24]  =  15'b001111110100111;     //24pi/512
   sin[25]  =  15'b111101100011100;     //25pi/512
   cos[25]  =  15'b001111110011111;     //25pi/512
   sin[26]  =  15'b111101011101011;     //26pi/512
   cos[26]  =  15'b001111110010111;     //26pi/512
   sin[27]  =  15'b111101010111001;     //27pi/512
   cos[27]  =  15'b001111110001111;     //27pi/512
   sin[28]  =  15'b111101010000111;     //28pi/512
   cos[28]  =  15'b001111110000111;     //28pi/512
   sin[29]  =  15'b111101001010110;     //29pi/512
   cos[29]  =  15'b001111101111110;     //29pi/512
   sin[30]  =  15'b111101000100101;     //30pi/512
   cos[30]  =  15'b001111101110101;     //30pi/512
   sin[31]  =  15'b111100111110011;     //31pi/512
   cos[31]  =  15'b001111101101100;     //31pi/512
   sin[32]  =  15'b111100111000010;     //32pi/512
   cos[32]  =  15'b001111101100010;     //32pi/512
   sin[33]  =  15'b111100110010001;     //33pi/512
   cos[33]  =  15'b001111101011000;     //33pi/512
   sin[34]  =  15'b111100101011111;     //34pi/512
   cos[34]  =  15'b001111101001110;     //34pi/512
   sin[35]  =  15'b111100100101110;     //35pi/512
   cos[35]  =  15'b001111101000011;     //35pi/512
   sin[36]  =  15'b111100011111101;     //36pi/512
   cos[36]  =  15'b001111100111000;     //36pi/512
   sin[37]  =  15'b111100011001100;     //37pi/512
   cos[37]  =  15'b001111100101101;     //37pi/512
   sin[38]  =  15'b111100010011011;     //38pi/512
   cos[38]  =  15'b001111100100010;     //38pi/512
   sin[39]  =  15'b111100001101010;     //39pi/512
   cos[39]  =  15'b001111100010110;     //39pi/512
   sin[40]  =  15'b111100000111010;     //40pi/512
   cos[40]  =  15'b001111100001010;     //40pi/512
   sin[41]  =  15'b111100000001001;     //41pi/512
   cos[41]  =  15'b001111011111110;     //41pi/512
   sin[42]  =  15'b111011111011000;     //42pi/512
   cos[42]  =  15'b001111011110001;     //42pi/512
   sin[43]  =  15'b111011110101000;     //43pi/512
   cos[43]  =  15'b001111011100100;     //43pi/512
   sin[44]  =  15'b111011101110111;     //44pi/512
   cos[44]  =  15'b001111011010111;     //44pi/512
   sin[45]  =  15'b111011101000111;     //45pi/512
   cos[45]  =  15'b001111011001001;     //45pi/512
   sin[46]  =  15'b111011100010110;     //46pi/512
   cos[46]  =  15'b001111010111011;     //46pi/512
   sin[47]  =  15'b111011011100110;     //47pi/512
   cos[47]  =  15'b001111010101101;     //47pi/512
   sin[48]  =  15'b111011010110110;     //48pi/512
   cos[48]  =  15'b001111010011111;     //48pi/512
   sin[49]  =  15'b111011010000110;     //49pi/512
   cos[49]  =  15'b001111010010000;     //49pi/512
   sin[50]  =  15'b111011001010110;     //50pi/512
   cos[50]  =  15'b001111010000001;     //50pi/512
   sin[51]  =  15'b111011000100110;     //51pi/512
   cos[51]  =  15'b001111001110010;     //51pi/512
   sin[52]  =  15'b111010111110110;     //52pi/512
   cos[52]  =  15'b001111001100010;     //52pi/512
   sin[53]  =  15'b111010111000111;     //53pi/512
   cos[53]  =  15'b001111001010010;     //53pi/512
   sin[54]  =  15'b111010110010111;     //54pi/512
   cos[54]  =  15'b001111001000010;     //54pi/512
   sin[55]  =  15'b111010101101000;     //55pi/512
   cos[55]  =  15'b001111000110001;     //55pi/512
   sin[56]  =  15'b111010100111000;     //56pi/512
   cos[56]  =  15'b001111000100001;     //56pi/512
   sin[57]  =  15'b111010100001001;     //57pi/512
   cos[57]  =  15'b001111000010000;     //57pi/512
   sin[58]  =  15'b111010011011010;     //58pi/512
   cos[58]  =  15'b001110111111110;     //58pi/512
   sin[59]  =  15'b111010010101011;     //59pi/512
   cos[59]  =  15'b001110111101101;     //59pi/512
   sin[60]  =  15'b111010001111100;     //60pi/512
   cos[60]  =  15'b001110111011011;     //60pi/512
   sin[61]  =  15'b111010001001101;     //61pi/512
   cos[61]  =  15'b001110111001000;     //61pi/512
   sin[62]  =  15'b111010000011110;     //62pi/512
   cos[62]  =  15'b001110110110110;     //62pi/512
   sin[63]  =  15'b111001111110000;     //63pi/512
   cos[63]  =  15'b001110110100011;     //63pi/512
   sin[64]  =  15'b111001111000001;     //64pi/512
   cos[64]  =  15'b001110110010000;     //64pi/512
   sin[65]  =  15'b111001110010011;     //65pi/512
   cos[65]  =  15'b001110101111101;     //65pi/512
   sin[66]  =  15'b111001101100100;     //66pi/512
   cos[66]  =  15'b001110101101001;     //66pi/512
   sin[67]  =  15'b111001100110110;     //67pi/512
   cos[67]  =  15'b001110101010101;     //67pi/512
   sin[68]  =  15'b111001100001000;     //68pi/512
   cos[68]  =  15'b001110101000001;     //68pi/512
   sin[69]  =  15'b111001011011010;     //69pi/512
   cos[69]  =  15'b001110100101100;     //69pi/512
   sin[70]  =  15'b111001010101101;     //70pi/512
   cos[70]  =  15'b001110100010111;     //70pi/512
   sin[71]  =  15'b111001001111111;     //71pi/512
   cos[71]  =  15'b001110100000010;     //71pi/512
   sin[72]  =  15'b111001001010001;     //72pi/512
   cos[72]  =  15'b001110011101101;     //72pi/512
   sin[73]  =  15'b111001000100100;     //73pi/512
   cos[73]  =  15'b001110011010111;     //73pi/512
   sin[74]  =  15'b111000111110111;     //74pi/512
   cos[74]  =  15'b001110011000001;     //74pi/512
   sin[75]  =  15'b111000111001010;     //75pi/512
   cos[75]  =  15'b001110010101011;     //75pi/512
   sin[76]  =  15'b111000110011101;     //76pi/512
   cos[76]  =  15'b001110010010101;     //76pi/512
   sin[77]  =  15'b111000101110000;     //77pi/512
   cos[77]  =  15'b001110001111110;     //77pi/512
   sin[78]  =  15'b111000101000011;     //78pi/512
   cos[78]  =  15'b001110001100111;     //78pi/512
   sin[79]  =  15'b111000100010111;     //79pi/512
   cos[79]  =  15'b001110001010000;     //79pi/512
   sin[80]  =  15'b111000011101010;     //80pi/512
   cos[80]  =  15'b001110000111000;     //80pi/512
   sin[81]  =  15'b111000010111110;     //81pi/512
   cos[81]  =  15'b001110000100000;     //81pi/512
   sin[82]  =  15'b111000010010010;     //82pi/512
   cos[82]  =  15'b001110000001000;     //82pi/512
   sin[83]  =  15'b111000001100110;     //83pi/512
   cos[83]  =  15'b001101111110000;     //83pi/512
   sin[84]  =  15'b111000000111010;     //84pi/512
   cos[84]  =  15'b001101111010111;     //84pi/512
   sin[85]  =  15'b111000000001111;     //85pi/512
   cos[85]  =  15'b001101110111110;     //85pi/512
   sin[86]  =  15'b110111111100011;     //86pi/512
   cos[86]  =  15'b001101110100101;     //86pi/512
   sin[87]  =  15'b110111110111000;     //87pi/512
   cos[87]  =  15'b001101110001100;     //87pi/512
   sin[88]  =  15'b110111110001100;     //88pi/512
   cos[88]  =  15'b001101101110010;     //88pi/512
   sin[89]  =  15'b110111101100001;     //89pi/512
   cos[89]  =  15'b001101101011000;     //89pi/512
   sin[90]  =  15'b110111100110111;     //90pi/512
   cos[90]  =  15'b001101100111110;     //90pi/512
   sin[91]  =  15'b110111100001100;     //91pi/512
   cos[91]  =  15'b001101100100011;     //91pi/512
   sin[92]  =  15'b110111011100001;     //92pi/512
   cos[92]  =  15'b001101100001001;     //92pi/512
   sin[93]  =  15'b110111010110111;     //93pi/512
   cos[93]  =  15'b001101011101110;     //93pi/512
   sin[94]  =  15'b110111010001101;     //94pi/512
   cos[94]  =  15'b001101011010010;     //94pi/512
   sin[95]  =  15'b110111001100011;     //95pi/512
   cos[95]  =  15'b001101010110111;     //95pi/512
   sin[96]  =  15'b110111000111001;     //96pi/512
   cos[96]  =  15'b001101010011011;     //96pi/512
   sin[97]  =  15'b110111000001111;     //97pi/512
   cos[97]  =  15'b001101001111111;     //97pi/512
   sin[98]  =  15'b110110111100110;     //98pi/512
   cos[98]  =  15'b001101001100011;     //98pi/512
   sin[99]  =  15'b110110110111100;     //99pi/512
   cos[99]  =  15'b001101001000110;     //99pi/512
   sin[100]  =  15'b110110110010011;     //100pi/512
   cos[100]  =  15'b001101000101001;     //100pi/512
   sin[101]  =  15'b110110101101010;     //101pi/512
   cos[101]  =  15'b001101000001100;     //101pi/512
   sin[102]  =  15'b110110101000001;     //102pi/512
   cos[102]  =  15'b001100111101111;     //102pi/512
   sin[103]  =  15'b110110100011000;     //103pi/512
   cos[103]  =  15'b001100111010001;     //103pi/512
   sin[104]  =  15'b110110011110000;     //104pi/512
   cos[104]  =  15'b001100110110011;     //104pi/512
   sin[105]  =  15'b110110011001000;     //105pi/512
   cos[105]  =  15'b001100110010101;     //105pi/512
   sin[106]  =  15'b110110010100000;     //106pi/512
   cos[106]  =  15'b001100101110111;     //106pi/512
   sin[107]  =  15'b110110001111000;     //107pi/512
   cos[107]  =  15'b001100101011000;     //107pi/512
   sin[108]  =  15'b110110001010000;     //108pi/512
   cos[108]  =  15'b001100100111010;     //108pi/512
   sin[109]  =  15'b110110000101000;     //109pi/512
   cos[109]  =  15'b001100100011011;     //109pi/512
   sin[110]  =  15'b110110000000001;     //110pi/512
   cos[110]  =  15'b001100011111011;     //110pi/512
   sin[111]  =  15'b110101111011010;     //111pi/512
   cos[111]  =  15'b001100011011100;     //111pi/512
   sin[112]  =  15'b110101110110011;     //112pi/512
   cos[112]  =  15'b001100010111100;     //112pi/512
   sin[113]  =  15'b110101110001100;     //113pi/512
   cos[113]  =  15'b001100010011100;     //113pi/512
   sin[114]  =  15'b110101101100110;     //114pi/512
   cos[114]  =  15'b001100001111100;     //114pi/512
   sin[115]  =  15'b110101100111111;     //115pi/512
   cos[115]  =  15'b001100001011011;     //115pi/512
   sin[116]  =  15'b110101100011001;     //116pi/512
   cos[116]  =  15'b001100000111011;     //116pi/512
   sin[117]  =  15'b110101011110011;     //117pi/512
   cos[117]  =  15'b001100000011010;     //117pi/512
   sin[118]  =  15'b110101011001101;     //118pi/512
   cos[118]  =  15'b001011111111000;     //118pi/512
   sin[119]  =  15'b110101010101000;     //119pi/512
   cos[119]  =  15'b001011111010111;     //119pi/512
   sin[120]  =  15'b110101010000011;     //120pi/512
   cos[120]  =  15'b001011110110101;     //120pi/512
   sin[121]  =  15'b110101001011101;     //121pi/512
   cos[121]  =  15'b001011110010100;     //121pi/512
   sin[122]  =  15'b110101000111001;     //122pi/512
   cos[122]  =  15'b001011101110001;     //122pi/512
   sin[123]  =  15'b110101000010100;     //123pi/512
   cos[123]  =  15'b001011101001111;     //123pi/512
   sin[124]  =  15'b110100111101111;     //124pi/512
   cos[124]  =  15'b001011100101101;     //124pi/512
   sin[125]  =  15'b110100111001011;     //125pi/512
   cos[125]  =  15'b001011100001010;     //125pi/512
   sin[126]  =  15'b110100110100111;     //126pi/512
   cos[126]  =  15'b001011011100111;     //126pi/512
   sin[127]  =  15'b110100110000011;     //127pi/512
   cos[127]  =  15'b001011011000100;     //127pi/512
   sin[128]  =  15'b110100101011111;     //128pi/512
   cos[128]  =  15'b001011010100000;     //128pi/512
   sin[129]  =  15'b110100100111100;     //129pi/512
   cos[129]  =  15'b001011001111100;     //129pi/512
   sin[130]  =  15'b110100100011001;     //130pi/512
   cos[130]  =  15'b001011001011001;     //130pi/512
   sin[131]  =  15'b110100011110110;     //131pi/512
   cos[131]  =  15'b001011000110101;     //131pi/512
   sin[132]  =  15'b110100011010011;     //132pi/512
   cos[132]  =  15'b001011000010000;     //132pi/512
   sin[133]  =  15'b110100010110000;     //133pi/512
   cos[133]  =  15'b001010111101100;     //133pi/512
   sin[134]  =  15'b110100010001110;     //134pi/512
   cos[134]  =  15'b001010111000111;     //134pi/512
   sin[135]  =  15'b110100001101100;     //135pi/512
   cos[135]  =  15'b001010110100010;     //135pi/512
   sin[136]  =  15'b110100001001010;     //136pi/512
   cos[136]  =  15'b001010101111101;     //136pi/512
   sin[137]  =  15'b110100000101000;     //137pi/512
   cos[137]  =  15'b001010101011000;     //137pi/512
   sin[138]  =  15'b110100000000111;     //138pi/512
   cos[138]  =  15'b001010100110010;     //138pi/512
   sin[139]  =  15'b110011111100110;     //139pi/512
   cos[139]  =  15'b001010100001100;     //139pi/512
   sin[140]  =  15'b110011111000101;     //140pi/512
   cos[140]  =  15'b001010011100110;     //140pi/512
   sin[141]  =  15'b110011110100100;     //141pi/512
   cos[141]  =  15'b001010011000000;     //141pi/512
   sin[142]  =  15'b110011110000100;     //142pi/512
   cos[142]  =  15'b001010010011010;     //142pi/512
   sin[143]  =  15'b110011101100100;     //143pi/512
   cos[143]  =  15'b001010001110011;     //143pi/512
   sin[144]  =  15'b110011101000011;     //144pi/512
   cos[144]  =  15'b001010001001100;     //144pi/512
   sin[145]  =  15'b110011100100100;     //145pi/512
   cos[145]  =  15'b001010000100101;     //145pi/512
   sin[146]  =  15'b110011100000100;     //146pi/512
   cos[146]  =  15'b001001111111110;     //146pi/512
   sin[147]  =  15'b110011011100101;     //147pi/512
   cos[147]  =  15'b001001111010111;     //147pi/512
   sin[148]  =  15'b110011011000110;     //148pi/512
   cos[148]  =  15'b001001110101111;     //148pi/512
   sin[149]  =  15'b110011010100111;     //149pi/512
   cos[149]  =  15'b001001110001000;     //149pi/512
   sin[150]  =  15'b110011010001001;     //150pi/512
   cos[150]  =  15'b001001101100000;     //150pi/512
   sin[151]  =  15'b110011001101010;     //151pi/512
   cos[151]  =  15'b001001100111000;     //151pi/512
   sin[152]  =  15'b110011001001100;     //152pi/512
   cos[152]  =  15'b001001100001111;     //152pi/512
   sin[153]  =  15'b110011000101110;     //153pi/512
   cos[153]  =  15'b001001011100111;     //153pi/512
   sin[154]  =  15'b110011000010001;     //154pi/512
   cos[154]  =  15'b001001010111110;     //154pi/512
   sin[155]  =  15'b110010111110011;     //155pi/512
   cos[155]  =  15'b001001010010110;     //155pi/512
   sin[156]  =  15'b110010111010110;     //156pi/512
   cos[156]  =  15'b001001001101101;     //156pi/512
   sin[157]  =  15'b110010110111010;     //157pi/512
   cos[157]  =  15'b001001001000011;     //157pi/512
   sin[158]  =  15'b110010110011101;     //158pi/512
   cos[158]  =  15'b001001000011010;     //158pi/512
   sin[159]  =  15'b110010110000001;     //159pi/512
   cos[159]  =  15'b001000111110000;     //159pi/512
   sin[160]  =  15'b110010101100101;     //160pi/512
   cos[160]  =  15'b001000111000111;     //160pi/512
   sin[161]  =  15'b110010101001001;     //161pi/512
   cos[161]  =  15'b001000110011101;     //161pi/512
   sin[162]  =  15'b110010100101101;     //162pi/512
   cos[162]  =  15'b001000101110011;     //162pi/512
   sin[163]  =  15'b110010100010010;     //163pi/512
   cos[163]  =  15'b001000101001001;     //163pi/512
   sin[164]  =  15'b110010011110111;     //164pi/512
   cos[164]  =  15'b001000100011110;     //164pi/512
   sin[165]  =  15'b110010011011100;     //165pi/512
   cos[165]  =  15'b001000011110100;     //165pi/512
   sin[166]  =  15'b110010011000010;     //166pi/512
   cos[166]  =  15'b001000011001001;     //166pi/512
   sin[167]  =  15'b110010010100111;     //167pi/512
   cos[167]  =  15'b001000010011110;     //167pi/512
   sin[168]  =  15'b110010010001101;     //168pi/512
   cos[168]  =  15'b001000001110011;     //168pi/512
   sin[169]  =  15'b110010001110100;     //169pi/512
   cos[169]  =  15'b001000001001000;     //169pi/512
   sin[170]  =  15'b110010001011010;     //170pi/512
   cos[170]  =  15'b001000000011100;     //170pi/512
   sin[171]  =  15'b110010001000001;     //171pi/512
   cos[171]  =  15'b000111111110001;     //171pi/512
   sin[172]  =  15'b110010000101000;     //172pi/512
   cos[172]  =  15'b000111111000101;     //172pi/512
   sin[173]  =  15'b110010000010000;     //173pi/512
   cos[173]  =  15'b000111110011010;     //173pi/512
   sin[174]  =  15'b110001111110111;     //174pi/512
   cos[174]  =  15'b000111101101110;     //174pi/512
   sin[175]  =  15'b110001111011111;     //175pi/512
   cos[175]  =  15'b000111101000001;     //175pi/512
   sin[176]  =  15'b110001111000111;     //176pi/512
   cos[176]  =  15'b000111100010101;     //176pi/512
   sin[177]  =  15'b110001110110000;     //177pi/512
   cos[177]  =  15'b000111011101001;     //177pi/512
   sin[178]  =  15'b110001110011000;     //178pi/512
   cos[178]  =  15'b000111010111100;     //178pi/512
   sin[179]  =  15'b110001110000001;     //179pi/512
   cos[179]  =  15'b000111010010000;     //179pi/512
   sin[180]  =  15'b110001101101011;     //180pi/512
   cos[180]  =  15'b000111001100011;     //180pi/512
   sin[181]  =  15'b110001101010100;     //181pi/512
   cos[181]  =  15'b000111000110110;     //181pi/512
   sin[182]  =  15'b110001100111110;     //182pi/512
   cos[182]  =  15'b000111000001001;     //182pi/512
   sin[183]  =  15'b110001100101000;     //183pi/512
   cos[183]  =  15'b000110111011011;     //183pi/512
   sin[184]  =  15'b110001100010011;     //184pi/512
   cos[184]  =  15'b000110110101110;     //184pi/512
   sin[185]  =  15'b110001011111101;     //185pi/512
   cos[185]  =  15'b000110110000001;     //185pi/512
   sin[186]  =  15'b110001011101000;     //186pi/512
   cos[186]  =  15'b000110101010011;     //186pi/512
   sin[187]  =  15'b110001011010011;     //187pi/512
   cos[187]  =  15'b000110100100101;     //187pi/512
   sin[188]  =  15'b110001010111111;     //188pi/512
   cos[188]  =  15'b000110011110111;     //188pi/512
   sin[189]  =  15'b110001010101011;     //189pi/512
   cos[189]  =  15'b000110011001001;     //189pi/512
   sin[190]  =  15'b110001010010111;     //190pi/512
   cos[190]  =  15'b000110010011011;     //190pi/512
   sin[191]  =  15'b110001010000011;     //191pi/512
   cos[191]  =  15'b000110001101101;     //191pi/512
   sin[192]  =  15'b110001001110000;     //192pi/512
   cos[192]  =  15'b000110000111110;     //192pi/512
   sin[193]  =  15'b110001001011100;     //193pi/512
   cos[193]  =  15'b000110000010000;     //193pi/512
   sin[194]  =  15'b110001001001010;     //194pi/512
   cos[194]  =  15'b000101111100001;     //194pi/512
   sin[195]  =  15'b110001000110111;     //195pi/512
   cos[195]  =  15'b000101110110011;     //195pi/512
   sin[196]  =  15'b110001000100101;     //196pi/512
   cos[196]  =  15'b000101110000100;     //196pi/512
   sin[197]  =  15'b110001000010011;     //197pi/512
   cos[197]  =  15'b000101101010101;     //197pi/512
   sin[198]  =  15'b110001000000001;     //198pi/512
   cos[198]  =  15'b000101100100110;     //198pi/512
   sin[199]  =  15'b110000111110000;     //199pi/512
   cos[199]  =  15'b000101011110111;     //199pi/512
   sin[200]  =  15'b110000111011111;     //200pi/512
   cos[200]  =  15'b000101011000111;     //200pi/512
   sin[201]  =  15'b110000111001110;     //201pi/512
   cos[201]  =  15'b000101010011000;     //201pi/512
   sin[202]  =  15'b110000110111110;     //202pi/512
   cos[202]  =  15'b000101001101000;     //202pi/512
   sin[203]  =  15'b110000110101101;     //203pi/512
   cos[203]  =  15'b000101000111001;     //203pi/512
   sin[204]  =  15'b110000110011101;     //204pi/512
   cos[204]  =  15'b000101000001001;     //204pi/512
   sin[205]  =  15'b110000110001110;     //205pi/512
   cos[205]  =  15'b000100111011001;     //205pi/512
   sin[206]  =  15'b110000101111111;     //206pi/512
   cos[206]  =  15'b000100110101010;     //206pi/512
   sin[207]  =  15'b110000101101111;     //207pi/512
   cos[207]  =  15'b000100101111010;     //207pi/512
   sin[208]  =  15'b110000101100001;     //208pi/512
   cos[208]  =  15'b000100101001010;     //208pi/512
   sin[209]  =  15'b110000101010010;     //209pi/512
   cos[209]  =  15'b000100100011001;     //209pi/512
   sin[210]  =  15'b110000101000100;     //210pi/512
   cos[210]  =  15'b000100011101001;     //210pi/512
   sin[211]  =  15'b110000100110110;     //211pi/512
   cos[211]  =  15'b000100010111001;     //211pi/512
   sin[212]  =  15'b110000100101001;     //212pi/512
   cos[212]  =  15'b000100010001000;     //212pi/512
   sin[213]  =  15'b110000100011011;     //213pi/512
   cos[213]  =  15'b000100001011000;     //213pi/512
   sin[214]  =  15'b110000100001111;     //214pi/512
   cos[214]  =  15'b000100000100111;     //214pi/512
   sin[215]  =  15'b110000100000010;     //215pi/512
   cos[215]  =  15'b000011111110111;     //215pi/512
   sin[216]  =  15'b110000011110110;     //216pi/512
   cos[216]  =  15'b000011111000110;     //216pi/512
   sin[217]  =  15'b110000011101001;     //217pi/512
   cos[217]  =  15'b000011110010101;     //217pi/512
   sin[218]  =  15'b110000011011110;     //218pi/512
   cos[218]  =  15'b000011101100100;     //218pi/512
   sin[219]  =  15'b110000011010010;     //219pi/512
   cos[219]  =  15'b000011100110011;     //219pi/512
   sin[220]  =  15'b110000011000111;     //220pi/512
   cos[220]  =  15'b000011100000010;     //220pi/512
   sin[221]  =  15'b110000010111100;     //221pi/512
   cos[221]  =  15'b000011011010001;     //221pi/512
   sin[222]  =  15'b110000010110010;     //222pi/512
   cos[222]  =  15'b000011010100000;     //222pi/512
   sin[223]  =  15'b110000010100111;     //223pi/512
   cos[223]  =  15'b000011001101111;     //223pi/512
   sin[224]  =  15'b110000010011101;     //224pi/512
   cos[224]  =  15'b000011000111110;     //224pi/512
   sin[225]  =  15'b110000010010100;     //225pi/512
   cos[225]  =  15'b000011000001100;     //225pi/512
   sin[226]  =  15'b110000010001010;     //226pi/512
   cos[226]  =  15'b000010111011011;     //226pi/512
   sin[227]  =  15'b110000010000001;     //227pi/512
   cos[227]  =  15'b000010110101010;     //227pi/512
   sin[228]  =  15'b110000001111001;     //228pi/512
   cos[228]  =  15'b000010101111000;     //228pi/512
   sin[229]  =  15'b110000001110000;     //229pi/512
   cos[229]  =  15'b000010101000110;     //229pi/512
   sin[230]  =  15'b110000001101000;     //230pi/512
   cos[230]  =  15'b000010100010101;     //230pi/512
   sin[231]  =  15'b110000001100000;     //231pi/512
   cos[231]  =  15'b000010011100011;     //231pi/512
   sin[232]  =  15'b110000001011001;     //232pi/512
   cos[232]  =  15'b000010010110010;     //232pi/512
   sin[233]  =  15'b110000001010001;     //233pi/512
   cos[233]  =  15'b000010010000000;     //233pi/512
   sin[234]  =  15'b110000001001011;     //234pi/512
   cos[234]  =  15'b000010001001110;     //234pi/512
   sin[235]  =  15'b110000001000100;     //235pi/512
   cos[235]  =  15'b000010000011100;     //235pi/512
   sin[236]  =  15'b110000000111110;     //236pi/512
   cos[236]  =  15'b000001111101010;     //236pi/512
   sin[237]  =  15'b110000000111000;     //237pi/512
   cos[237]  =  15'b000001110111000;     //237pi/512
   sin[238]  =  15'b110000000110010;     //238pi/512
   cos[238]  =  15'b000001110000110;     //238pi/512
   sin[239]  =  15'b110000000101101;     //239pi/512
   cos[239]  =  15'b000001101010100;     //239pi/512
   sin[240]  =  15'b110000000100111;     //240pi/512
   cos[240]  =  15'b000001100100010;     //240pi/512
   sin[241]  =  15'b110000000100011;     //241pi/512
   cos[241]  =  15'b000001011110000;     //241pi/512
   sin[242]  =  15'b110000000011110;     //242pi/512
   cos[242]  =  15'b000001010111110;     //242pi/512
   sin[243]  =  15'b110000000011010;     //243pi/512
   cos[243]  =  15'b000001010001100;     //243pi/512
   sin[244]  =  15'b110000000010110;     //244pi/512
   cos[244]  =  15'b000001001011010;     //244pi/512
   sin[245]  =  15'b110000000010011;     //245pi/512
   cos[245]  =  15'b000001000101000;     //245pi/512
   sin[246]  =  15'b110000000001111;     //246pi/512
   cos[246]  =  15'b000000111110110;     //246pi/512
   sin[247]  =  15'b110000000001100;     //247pi/512
   cos[247]  =  15'b000000111000100;     //247pi/512
   sin[248]  =  15'b110000000001010;     //248pi/512
   cos[248]  =  15'b000000110010001;     //248pi/512
   sin[249]  =  15'b110000000001000;     //249pi/512
   cos[249]  =  15'b000000101011111;     //249pi/512
   sin[250]  =  15'b110000000000110;     //250pi/512
   cos[250]  =  15'b000000100101101;     //250pi/512
   sin[251]  =  15'b110000000000100;     //251pi/512
   cos[251]  =  15'b000000011111011;     //251pi/512
   sin[252]  =  15'b110000000000010;     //252pi/512
   cos[252]  =  15'b000000011001001;     //252pi/512
   sin[253]  =  15'b110000000000001;     //253pi/512
   cos[253]  =  15'b000000010010110;     //253pi/512
   sin[254]  =  15'b110000000000001;     //254pi/512
   cos[254]  =  15'b000000001100100;     //254pi/512
   sin[255]  =  15'b110000000000000;     //255pi/512
   cos[255]  =  15'b000000000110010;     //255pi/512
   sin[256]  =  15'b110000000000000;     //256pi/512
   cos[256]  =  15'b000000000000000;     //256pi/512
   sin[257]  =  15'b110000000000000;     //257pi/512
   cos[257]  =  15'b111111111001110;     //257pi/512
   sin[258]  =  15'b110000000000001;     //258pi/512
   cos[258]  =  15'b111111110011011;     //258pi/512
   sin[259]  =  15'b110000000000001;     //259pi/512
   cos[259]  =  15'b111111101101001;     //259pi/512
   sin[260]  =  15'b110000000000010;     //260pi/512
   cos[260]  =  15'b111111100110111;     //260pi/512
   sin[261]  =  15'b110000000000100;     //261pi/512
   cos[261]  =  15'b111111100000101;     //261pi/512
   sin[262]  =  15'b110000000000110;     //262pi/512
   cos[262]  =  15'b111111011010010;     //262pi/512
   sin[263]  =  15'b110000000001000;     //263pi/512
   cos[263]  =  15'b111111010100000;     //263pi/512
   sin[264]  =  15'b110000000001010;     //264pi/512
   cos[264]  =  15'b111111001101110;     //264pi/512
   sin[265]  =  15'b110000000001100;     //265pi/512
   cos[265]  =  15'b111111000111100;     //265pi/512
   sin[266]  =  15'b110000000001111;     //266pi/512
   cos[266]  =  15'b111111000001010;     //266pi/512
   sin[267]  =  15'b110000000010011;     //267pi/512
   cos[267]  =  15'b111110111010111;     //267pi/512
   sin[268]  =  15'b110000000010110;     //268pi/512
   cos[268]  =  15'b111110110100101;     //268pi/512
   sin[269]  =  15'b110000000011010;     //269pi/512
   cos[269]  =  15'b111110101110011;     //269pi/512
   sin[270]  =  15'b110000000011110;     //270pi/512
   cos[270]  =  15'b111110101000001;     //270pi/512
   sin[271]  =  15'b110000000100011;     //271pi/512
   cos[271]  =  15'b111110100001111;     //271pi/512
   sin[272]  =  15'b110000000100111;     //272pi/512
   cos[272]  =  15'b111110011011101;     //272pi/512
   sin[273]  =  15'b110000000101101;     //273pi/512
   cos[273]  =  15'b111110010101011;     //273pi/512
   sin[274]  =  15'b110000000110010;     //274pi/512
   cos[274]  =  15'b111110001111001;     //274pi/512
   sin[275]  =  15'b110000000111000;     //275pi/512
   cos[275]  =  15'b111110001000111;     //275pi/512
   sin[276]  =  15'b110000000111110;     //276pi/512
   cos[276]  =  15'b111110000010101;     //276pi/512
   sin[277]  =  15'b110000001000100;     //277pi/512
   cos[277]  =  15'b111101111100011;     //277pi/512
   sin[278]  =  15'b110000001001011;     //278pi/512
   cos[278]  =  15'b111101110110010;     //278pi/512
   sin[279]  =  15'b110000001010001;     //279pi/512
   cos[279]  =  15'b111101110000000;     //279pi/512
   sin[280]  =  15'b110000001011001;     //280pi/512
   cos[280]  =  15'b111101101001110;     //280pi/512
   sin[281]  =  15'b110000001100000;     //281pi/512
   cos[281]  =  15'b111101100011100;     //281pi/512
   sin[282]  =  15'b110000001101000;     //282pi/512
   cos[282]  =  15'b111101011101011;     //282pi/512
   sin[283]  =  15'b110000001110000;     //283pi/512
   cos[283]  =  15'b111101010111001;     //283pi/512
   sin[284]  =  15'b110000001111001;     //284pi/512
   cos[284]  =  15'b111101010000111;     //284pi/512
   sin[285]  =  15'b110000010000001;     //285pi/512
   cos[285]  =  15'b111101001010110;     //285pi/512
   sin[286]  =  15'b110000010001010;     //286pi/512
   cos[286]  =  15'b111101000100101;     //286pi/512
   sin[287]  =  15'b110000010010100;     //287pi/512
   cos[287]  =  15'b111100111110011;     //287pi/512
   sin[288]  =  15'b110000010011101;     //288pi/512
   cos[288]  =  15'b111100111000010;     //288pi/512
   sin[289]  =  15'b110000010100111;     //289pi/512
   cos[289]  =  15'b111100110010001;     //289pi/512
   sin[290]  =  15'b110000010110010;     //290pi/512
   cos[290]  =  15'b111100101011111;     //290pi/512
   sin[291]  =  15'b110000010111100;     //291pi/512
   cos[291]  =  15'b111100100101110;     //291pi/512
   sin[292]  =  15'b110000011000111;     //292pi/512
   cos[292]  =  15'b111100011111101;     //292pi/512
   sin[293]  =  15'b110000011010010;     //293pi/512
   cos[293]  =  15'b111100011001100;     //293pi/512
   sin[294]  =  15'b110000011011110;     //294pi/512
   cos[294]  =  15'b111100010011011;     //294pi/512
   sin[295]  =  15'b110000011101001;     //295pi/512
   cos[295]  =  15'b111100001101010;     //295pi/512
   sin[296]  =  15'b110000011110110;     //296pi/512
   cos[296]  =  15'b111100000111010;     //296pi/512
   sin[297]  =  15'b110000100000010;     //297pi/512
   cos[297]  =  15'b111100000001001;     //297pi/512
   sin[298]  =  15'b110000100001111;     //298pi/512
   cos[298]  =  15'b111011111011000;     //298pi/512
   sin[299]  =  15'b110000100011011;     //299pi/512
   cos[299]  =  15'b111011110101000;     //299pi/512
   sin[300]  =  15'b110000100101001;     //300pi/512
   cos[300]  =  15'b111011101110111;     //300pi/512
   sin[301]  =  15'b110000100110110;     //301pi/512
   cos[301]  =  15'b111011101000111;     //301pi/512
   sin[302]  =  15'b110000101000100;     //302pi/512
   cos[302]  =  15'b111011100010110;     //302pi/512
   sin[303]  =  15'b110000101010010;     //303pi/512
   cos[303]  =  15'b111011011100110;     //303pi/512
   sin[304]  =  15'b110000101100001;     //304pi/512
   cos[304]  =  15'b111011010110110;     //304pi/512
   sin[305]  =  15'b110000101101111;     //305pi/512
   cos[305]  =  15'b111011010000110;     //305pi/512
   sin[306]  =  15'b110000101111111;     //306pi/512
   cos[306]  =  15'b111011001010110;     //306pi/512
   sin[307]  =  15'b110000110001110;     //307pi/512
   cos[307]  =  15'b111011000100110;     //307pi/512
   sin[308]  =  15'b110000110011101;     //308pi/512
   cos[308]  =  15'b111010111110110;     //308pi/512
   sin[309]  =  15'b110000110101101;     //309pi/512
   cos[309]  =  15'b111010111000111;     //309pi/512
   sin[310]  =  15'b110000110111110;     //310pi/512
   cos[310]  =  15'b111010110010111;     //310pi/512
   sin[311]  =  15'b110000111001110;     //311pi/512
   cos[311]  =  15'b111010101101000;     //311pi/512
   sin[312]  =  15'b110000111011111;     //312pi/512
   cos[312]  =  15'b111010100111000;     //312pi/512
   sin[313]  =  15'b110000111110000;     //313pi/512
   cos[313]  =  15'b111010100001001;     //313pi/512
   sin[314]  =  15'b110001000000001;     //314pi/512
   cos[314]  =  15'b111010011011010;     //314pi/512
   sin[315]  =  15'b110001000010011;     //315pi/512
   cos[315]  =  15'b111010010101011;     //315pi/512
   sin[316]  =  15'b110001000100101;     //316pi/512
   cos[316]  =  15'b111010001111100;     //316pi/512
   sin[317]  =  15'b110001000110111;     //317pi/512
   cos[317]  =  15'b111010001001101;     //317pi/512
   sin[318]  =  15'b110001001001010;     //318pi/512
   cos[318]  =  15'b111010000011110;     //318pi/512
   sin[319]  =  15'b110001001011100;     //319pi/512
   cos[319]  =  15'b111001111110000;     //319pi/512
   sin[320]  =  15'b110001001110000;     //320pi/512
   cos[320]  =  15'b111001111000001;     //320pi/512
   sin[321]  =  15'b110001010000011;     //321pi/512
   cos[321]  =  15'b111001110010011;     //321pi/512
   sin[322]  =  15'b110001010010111;     //322pi/512
   cos[322]  =  15'b111001101100100;     //322pi/512
   sin[323]  =  15'b110001010101011;     //323pi/512
   cos[323]  =  15'b111001100110110;     //323pi/512
   sin[324]  =  15'b110001010111111;     //324pi/512
   cos[324]  =  15'b111001100001000;     //324pi/512
   sin[325]  =  15'b110001011010011;     //325pi/512
   cos[325]  =  15'b111001011011010;     //325pi/512
   sin[326]  =  15'b110001011101000;     //326pi/512
   cos[326]  =  15'b111001010101101;     //326pi/512
   sin[327]  =  15'b110001011111101;     //327pi/512
   cos[327]  =  15'b111001001111111;     //327pi/512
   sin[328]  =  15'b110001100010011;     //328pi/512
   cos[328]  =  15'b111001001010001;     //328pi/512
   sin[329]  =  15'b110001100101000;     //329pi/512
   cos[329]  =  15'b111001000100100;     //329pi/512
   sin[330]  =  15'b110001100111110;     //330pi/512
   cos[330]  =  15'b111000111110111;     //330pi/512
   sin[331]  =  15'b110001101010100;     //331pi/512
   cos[331]  =  15'b111000111001010;     //331pi/512
   sin[332]  =  15'b110001101101011;     //332pi/512
   cos[332]  =  15'b111000110011101;     //332pi/512
   sin[333]  =  15'b110001110000001;     //333pi/512
   cos[333]  =  15'b111000101110000;     //333pi/512
   sin[334]  =  15'b110001110011000;     //334pi/512
   cos[334]  =  15'b111000101000011;     //334pi/512
   sin[335]  =  15'b110001110110000;     //335pi/512
   cos[335]  =  15'b111000100010111;     //335pi/512
   sin[336]  =  15'b110001111000111;     //336pi/512
   cos[336]  =  15'b111000011101010;     //336pi/512
   sin[337]  =  15'b110001111011111;     //337pi/512
   cos[337]  =  15'b111000010111110;     //337pi/512
   sin[338]  =  15'b110001111110111;     //338pi/512
   cos[338]  =  15'b111000010010010;     //338pi/512
   sin[339]  =  15'b110010000010000;     //339pi/512
   cos[339]  =  15'b111000001100110;     //339pi/512
   sin[340]  =  15'b110010000101000;     //340pi/512
   cos[340]  =  15'b111000000111010;     //340pi/512
   sin[341]  =  15'b110010001000001;     //341pi/512
   cos[341]  =  15'b111000000001111;     //341pi/512
   sin[342]  =  15'b110010001011010;     //342pi/512
   cos[342]  =  15'b110111111100011;     //342pi/512
   sin[343]  =  15'b110010001110100;     //343pi/512
   cos[343]  =  15'b110111110111000;     //343pi/512
   sin[344]  =  15'b110010010001101;     //344pi/512
   cos[344]  =  15'b110111110001100;     //344pi/512
   sin[345]  =  15'b110010010100111;     //345pi/512
   cos[345]  =  15'b110111101100001;     //345pi/512
   sin[346]  =  15'b110010011000010;     //346pi/512
   cos[346]  =  15'b110111100110111;     //346pi/512
   sin[347]  =  15'b110010011011100;     //347pi/512
   cos[347]  =  15'b110111100001100;     //347pi/512
   sin[348]  =  15'b110010011110111;     //348pi/512
   cos[348]  =  15'b110111011100001;     //348pi/512
   sin[349]  =  15'b110010100010010;     //349pi/512
   cos[349]  =  15'b110111010110111;     //349pi/512
   sin[350]  =  15'b110010100101101;     //350pi/512
   cos[350]  =  15'b110111010001101;     //350pi/512
   sin[351]  =  15'b110010101001001;     //351pi/512
   cos[351]  =  15'b110111001100011;     //351pi/512
   sin[352]  =  15'b110010101100101;     //352pi/512
   cos[352]  =  15'b110111000111001;     //352pi/512
   sin[353]  =  15'b110010110000001;     //353pi/512
   cos[353]  =  15'b110111000001111;     //353pi/512
   sin[354]  =  15'b110010110011101;     //354pi/512
   cos[354]  =  15'b110110111100110;     //354pi/512
   sin[355]  =  15'b110010110111010;     //355pi/512
   cos[355]  =  15'b110110110111100;     //355pi/512
   sin[356]  =  15'b110010111010110;     //356pi/512
   cos[356]  =  15'b110110110010011;     //356pi/512
   sin[357]  =  15'b110010111110011;     //357pi/512
   cos[357]  =  15'b110110101101010;     //357pi/512
   sin[358]  =  15'b110011000010001;     //358pi/512
   cos[358]  =  15'b110110101000001;     //358pi/512
   sin[359]  =  15'b110011000101110;     //359pi/512
   cos[359]  =  15'b110110100011000;     //359pi/512
   sin[360]  =  15'b110011001001100;     //360pi/512
   cos[360]  =  15'b110110011110000;     //360pi/512
   sin[361]  =  15'b110011001101010;     //361pi/512
   cos[361]  =  15'b110110011001000;     //361pi/512
   sin[362]  =  15'b110011010001001;     //362pi/512
   cos[362]  =  15'b110110010100000;     //362pi/512
   sin[363]  =  15'b110011010100111;     //363pi/512
   cos[363]  =  15'b110110001111000;     //363pi/512
   sin[364]  =  15'b110011011000110;     //364pi/512
   cos[364]  =  15'b110110001010000;     //364pi/512
   sin[365]  =  15'b110011011100101;     //365pi/512
   cos[365]  =  15'b110110000101000;     //365pi/512
   sin[366]  =  15'b110011100000100;     //366pi/512
   cos[366]  =  15'b110110000000001;     //366pi/512
   sin[367]  =  15'b110011100100100;     //367pi/512
   cos[367]  =  15'b110101111011010;     //367pi/512
   sin[368]  =  15'b110011101000011;     //368pi/512
   cos[368]  =  15'b110101110110011;     //368pi/512
   sin[369]  =  15'b110011101100100;     //369pi/512
   cos[369]  =  15'b110101110001100;     //369pi/512
   sin[370]  =  15'b110011110000100;     //370pi/512
   cos[370]  =  15'b110101101100110;     //370pi/512
   sin[371]  =  15'b110011110100100;     //371pi/512
   cos[371]  =  15'b110101100111111;     //371pi/512
   sin[372]  =  15'b110011111000101;     //372pi/512
   cos[372]  =  15'b110101100011001;     //372pi/512
   sin[373]  =  15'b110011111100110;     //373pi/512
   cos[373]  =  15'b110101011110011;     //373pi/512
   sin[374]  =  15'b110100000000111;     //374pi/512
   cos[374]  =  15'b110101011001101;     //374pi/512
   sin[375]  =  15'b110100000101000;     //375pi/512
   cos[375]  =  15'b110101010101000;     //375pi/512
   sin[376]  =  15'b110100001001010;     //376pi/512
   cos[376]  =  15'b110101010000011;     //376pi/512
   sin[377]  =  15'b110100001101100;     //377pi/512
   cos[377]  =  15'b110101001011101;     //377pi/512
   sin[378]  =  15'b110100010001110;     //378pi/512
   cos[378]  =  15'b110101000111001;     //378pi/512
   sin[379]  =  15'b110100010110000;     //379pi/512
   cos[379]  =  15'b110101000010100;     //379pi/512
   sin[380]  =  15'b110100011010011;     //380pi/512
   cos[380]  =  15'b110100111101111;     //380pi/512
   sin[381]  =  15'b110100011110110;     //381pi/512
   cos[381]  =  15'b110100111001011;     //381pi/512
   sin[382]  =  15'b110100100011001;     //382pi/512
   cos[382]  =  15'b110100110100111;     //382pi/512
   sin[383]  =  15'b110100100111100;     //383pi/512
   cos[383]  =  15'b110100110000011;     //383pi/512
   sin[384]  =  15'b110100101011111;     //384pi/512
   cos[384]  =  15'b110100101011111;     //384pi/512
   sin[385]  =  15'b110100110000011;     //385pi/512
   cos[385]  =  15'b110100100111100;     //385pi/512
   sin[386]  =  15'b110100110100111;     //386pi/512
   cos[386]  =  15'b110100100011001;     //386pi/512
   sin[387]  =  15'b110100111001011;     //387pi/512
   cos[387]  =  15'b110100011110110;     //387pi/512
   sin[388]  =  15'b110100111101111;     //388pi/512
   cos[388]  =  15'b110100011010011;     //388pi/512
   sin[389]  =  15'b110101000010100;     //389pi/512
   cos[389]  =  15'b110100010110000;     //389pi/512
   sin[390]  =  15'b110101000111001;     //390pi/512
   cos[390]  =  15'b110100010001110;     //390pi/512
   sin[391]  =  15'b110101001011101;     //391pi/512
   cos[391]  =  15'b110100001101100;     //391pi/512
   sin[392]  =  15'b110101010000011;     //392pi/512
   cos[392]  =  15'b110100001001010;     //392pi/512
   sin[393]  =  15'b110101010101000;     //393pi/512
   cos[393]  =  15'b110100000101000;     //393pi/512
   sin[394]  =  15'b110101011001101;     //394pi/512
   cos[394]  =  15'b110100000000111;     //394pi/512
   sin[395]  =  15'b110101011110011;     //395pi/512
   cos[395]  =  15'b110011111100110;     //395pi/512
   sin[396]  =  15'b110101100011001;     //396pi/512
   cos[396]  =  15'b110011111000101;     //396pi/512
   sin[397]  =  15'b110101100111111;     //397pi/512
   cos[397]  =  15'b110011110100100;     //397pi/512
   sin[398]  =  15'b110101101100110;     //398pi/512
   cos[398]  =  15'b110011110000100;     //398pi/512
   sin[399]  =  15'b110101110001100;     //399pi/512
   cos[399]  =  15'b110011101100100;     //399pi/512
   sin[400]  =  15'b110101110110011;     //400pi/512
   cos[400]  =  15'b110011101000011;     //400pi/512
   sin[401]  =  15'b110101111011010;     //401pi/512
   cos[401]  =  15'b110011100100100;     //401pi/512
   sin[402]  =  15'b110110000000001;     //402pi/512
   cos[402]  =  15'b110011100000100;     //402pi/512
   sin[403]  =  15'b110110000101000;     //403pi/512
   cos[403]  =  15'b110011011100101;     //403pi/512
   sin[404]  =  15'b110110001010000;     //404pi/512
   cos[404]  =  15'b110011011000110;     //404pi/512
   sin[405]  =  15'b110110001111000;     //405pi/512
   cos[405]  =  15'b110011010100111;     //405pi/512
   sin[406]  =  15'b110110010100000;     //406pi/512
   cos[406]  =  15'b110011010001001;     //406pi/512
   sin[407]  =  15'b110110011001000;     //407pi/512
   cos[407]  =  15'b110011001101010;     //407pi/512
   sin[408]  =  15'b110110011110000;     //408pi/512
   cos[408]  =  15'b110011001001100;     //408pi/512
   sin[409]  =  15'b110110100011000;     //409pi/512
   cos[409]  =  15'b110011000101110;     //409pi/512
   sin[410]  =  15'b110110101000001;     //410pi/512
   cos[410]  =  15'b110011000010001;     //410pi/512
   sin[411]  =  15'b110110101101010;     //411pi/512
   cos[411]  =  15'b110010111110011;     //411pi/512
   sin[412]  =  15'b110110110010011;     //412pi/512
   cos[412]  =  15'b110010111010110;     //412pi/512
   sin[413]  =  15'b110110110111100;     //413pi/512
   cos[413]  =  15'b110010110111010;     //413pi/512
   sin[414]  =  15'b110110111100110;     //414pi/512
   cos[414]  =  15'b110010110011101;     //414pi/512
   sin[415]  =  15'b110111000001111;     //415pi/512
   cos[415]  =  15'b110010110000001;     //415pi/512
   sin[416]  =  15'b110111000111001;     //416pi/512
   cos[416]  =  15'b110010101100101;     //416pi/512
   sin[417]  =  15'b110111001100011;     //417pi/512
   cos[417]  =  15'b110010101001001;     //417pi/512
   sin[418]  =  15'b110111010001101;     //418pi/512
   cos[418]  =  15'b110010100101101;     //418pi/512
   sin[419]  =  15'b110111010110111;     //419pi/512
   cos[419]  =  15'b110010100010010;     //419pi/512
   sin[420]  =  15'b110111011100001;     //420pi/512
   cos[420]  =  15'b110010011110111;     //420pi/512
   sin[421]  =  15'b110111100001100;     //421pi/512
   cos[421]  =  15'b110010011011100;     //421pi/512
   sin[422]  =  15'b110111100110111;     //422pi/512
   cos[422]  =  15'b110010011000010;     //422pi/512
   sin[423]  =  15'b110111101100001;     //423pi/512
   cos[423]  =  15'b110010010100111;     //423pi/512
   sin[424]  =  15'b110111110001100;     //424pi/512
   cos[424]  =  15'b110010010001101;     //424pi/512
   sin[425]  =  15'b110111110111000;     //425pi/512
   cos[425]  =  15'b110010001110100;     //425pi/512
   sin[426]  =  15'b110111111100011;     //426pi/512
   cos[426]  =  15'b110010001011010;     //426pi/512
   sin[427]  =  15'b111000000001111;     //427pi/512
   cos[427]  =  15'b110010001000001;     //427pi/512
   sin[428]  =  15'b111000000111010;     //428pi/512
   cos[428]  =  15'b110010000101000;     //428pi/512
   sin[429]  =  15'b111000001100110;     //429pi/512
   cos[429]  =  15'b110010000010000;     //429pi/512
   sin[430]  =  15'b111000010010010;     //430pi/512
   cos[430]  =  15'b110001111110111;     //430pi/512
   sin[431]  =  15'b111000010111110;     //431pi/512
   cos[431]  =  15'b110001111011111;     //431pi/512
   sin[432]  =  15'b111000011101010;     //432pi/512
   cos[432]  =  15'b110001111000111;     //432pi/512
   sin[433]  =  15'b111000100010111;     //433pi/512
   cos[433]  =  15'b110001110110000;     //433pi/512
   sin[434]  =  15'b111000101000011;     //434pi/512
   cos[434]  =  15'b110001110011000;     //434pi/512
   sin[435]  =  15'b111000101110000;     //435pi/512
   cos[435]  =  15'b110001110000001;     //435pi/512
   sin[436]  =  15'b111000110011101;     //436pi/512
   cos[436]  =  15'b110001101101011;     //436pi/512
   sin[437]  =  15'b111000111001010;     //437pi/512
   cos[437]  =  15'b110001101010100;     //437pi/512
   sin[438]  =  15'b111000111110111;     //438pi/512
   cos[438]  =  15'b110001100111110;     //438pi/512
   sin[439]  =  15'b111001000100100;     //439pi/512
   cos[439]  =  15'b110001100101000;     //439pi/512
   sin[440]  =  15'b111001001010001;     //440pi/512
   cos[440]  =  15'b110001100010011;     //440pi/512
   sin[441]  =  15'b111001001111111;     //441pi/512
   cos[441]  =  15'b110001011111101;     //441pi/512
   sin[442]  =  15'b111001010101101;     //442pi/512
   cos[442]  =  15'b110001011101000;     //442pi/512
   sin[443]  =  15'b111001011011010;     //443pi/512
   cos[443]  =  15'b110001011010011;     //443pi/512
   sin[444]  =  15'b111001100001000;     //444pi/512
   cos[444]  =  15'b110001010111111;     //444pi/512
   sin[445]  =  15'b111001100110110;     //445pi/512
   cos[445]  =  15'b110001010101011;     //445pi/512
   sin[446]  =  15'b111001101100100;     //446pi/512
   cos[446]  =  15'b110001010010111;     //446pi/512
   sin[447]  =  15'b111001110010011;     //447pi/512
   cos[447]  =  15'b110001010000011;     //447pi/512
   sin[448]  =  15'b111001111000001;     //448pi/512
   cos[448]  =  15'b110001001110000;     //448pi/512
   sin[449]  =  15'b111001111110000;     //449pi/512
   cos[449]  =  15'b110001001011100;     //449pi/512
   sin[450]  =  15'b111010000011110;     //450pi/512
   cos[450]  =  15'b110001001001010;     //450pi/512
   sin[451]  =  15'b111010001001101;     //451pi/512
   cos[451]  =  15'b110001000110111;     //451pi/512
   sin[452]  =  15'b111010001111100;     //452pi/512
   cos[452]  =  15'b110001000100101;     //452pi/512
   sin[453]  =  15'b111010010101011;     //453pi/512
   cos[453]  =  15'b110001000010011;     //453pi/512
   sin[454]  =  15'b111010011011010;     //454pi/512
   cos[454]  =  15'b110001000000001;     //454pi/512
   sin[455]  =  15'b111010100001001;     //455pi/512
   cos[455]  =  15'b110000111110000;     //455pi/512
   sin[456]  =  15'b111010100111000;     //456pi/512
   cos[456]  =  15'b110000111011111;     //456pi/512
   sin[457]  =  15'b111010101101000;     //457pi/512
   cos[457]  =  15'b110000111001110;     //457pi/512
   sin[458]  =  15'b111010110010111;     //458pi/512
   cos[458]  =  15'b110000110111110;     //458pi/512
   sin[459]  =  15'b111010111000111;     //459pi/512
   cos[459]  =  15'b110000110101101;     //459pi/512
   sin[460]  =  15'b111010111110110;     //460pi/512
   cos[460]  =  15'b110000110011101;     //460pi/512
   sin[461]  =  15'b111011000100110;     //461pi/512
   cos[461]  =  15'b110000110001110;     //461pi/512
   sin[462]  =  15'b111011001010110;     //462pi/512
   cos[462]  =  15'b110000101111111;     //462pi/512
   sin[463]  =  15'b111011010000110;     //463pi/512
   cos[463]  =  15'b110000101101111;     //463pi/512
   sin[464]  =  15'b111011010110110;     //464pi/512
   cos[464]  =  15'b110000101100001;     //464pi/512
   sin[465]  =  15'b111011011100110;     //465pi/512
   cos[465]  =  15'b110000101010010;     //465pi/512
   sin[466]  =  15'b111011100010110;     //466pi/512
   cos[466]  =  15'b110000101000100;     //466pi/512
   sin[467]  =  15'b111011101000111;     //467pi/512
   cos[467]  =  15'b110000100110110;     //467pi/512
   sin[468]  =  15'b111011101110111;     //468pi/512
   cos[468]  =  15'b110000100101001;     //468pi/512
   sin[469]  =  15'b111011110101000;     //469pi/512
   cos[469]  =  15'b110000100011011;     //469pi/512
   sin[470]  =  15'b111011111011000;     //470pi/512
   cos[470]  =  15'b110000100001111;     //470pi/512
   sin[471]  =  15'b111100000001001;     //471pi/512
   cos[471]  =  15'b110000100000010;     //471pi/512
   sin[472]  =  15'b111100000111010;     //472pi/512
   cos[472]  =  15'b110000011110110;     //472pi/512
   sin[473]  =  15'b111100001101010;     //473pi/512
   cos[473]  =  15'b110000011101001;     //473pi/512
   sin[474]  =  15'b111100010011011;     //474pi/512
   cos[474]  =  15'b110000011011110;     //474pi/512
   sin[475]  =  15'b111100011001100;     //475pi/512
   cos[475]  =  15'b110000011010010;     //475pi/512
   sin[476]  =  15'b111100011111101;     //476pi/512
   cos[476]  =  15'b110000011000111;     //476pi/512
   sin[477]  =  15'b111100100101110;     //477pi/512
   cos[477]  =  15'b110000010111100;     //477pi/512
   sin[478]  =  15'b111100101011111;     //478pi/512
   cos[478]  =  15'b110000010110010;     //478pi/512
   sin[479]  =  15'b111100110010001;     //479pi/512
   cos[479]  =  15'b110000010100111;     //479pi/512
   sin[480]  =  15'b111100111000010;     //480pi/512
   cos[480]  =  15'b110000010011101;     //480pi/512
   sin[481]  =  15'b111100111110011;     //481pi/512
   cos[481]  =  15'b110000010010100;     //481pi/512
   sin[482]  =  15'b111101000100101;     //482pi/512
   cos[482]  =  15'b110000010001010;     //482pi/512
   sin[483]  =  15'b111101001010110;     //483pi/512
   cos[483]  =  15'b110000010000001;     //483pi/512
   sin[484]  =  15'b111101010000111;     //484pi/512
   cos[484]  =  15'b110000001111001;     //484pi/512
   sin[485]  =  15'b111101010111001;     //485pi/512
   cos[485]  =  15'b110000001110000;     //485pi/512
   sin[486]  =  15'b111101011101011;     //486pi/512
   cos[486]  =  15'b110000001101000;     //486pi/512
   sin[487]  =  15'b111101100011100;     //487pi/512
   cos[487]  =  15'b110000001100000;     //487pi/512
   sin[488]  =  15'b111101101001110;     //488pi/512
   cos[488]  =  15'b110000001011001;     //488pi/512
   sin[489]  =  15'b111101110000000;     //489pi/512
   cos[489]  =  15'b110000001010001;     //489pi/512
   sin[490]  =  15'b111101110110010;     //490pi/512
   cos[490]  =  15'b110000001001011;     //490pi/512
   sin[491]  =  15'b111101111100011;     //491pi/512
   cos[491]  =  15'b110000001000100;     //491pi/512
   sin[492]  =  15'b111110000010101;     //492pi/512
   cos[492]  =  15'b110000000111110;     //492pi/512
   sin[493]  =  15'b111110001000111;     //493pi/512
   cos[493]  =  15'b110000000111000;     //493pi/512
   sin[494]  =  15'b111110001111001;     //494pi/512
   cos[494]  =  15'b110000000110010;     //494pi/512
   sin[495]  =  15'b111110010101011;     //495pi/512
   cos[495]  =  15'b110000000101101;     //495pi/512
   sin[496]  =  15'b111110011011101;     //496pi/512
   cos[496]  =  15'b110000000100111;     //496pi/512
   sin[497]  =  15'b111110100001111;     //497pi/512
   cos[497]  =  15'b110000000100011;     //497pi/512
   sin[498]  =  15'b111110101000001;     //498pi/512
   cos[498]  =  15'b110000000011110;     //498pi/512
   sin[499]  =  15'b111110101110011;     //499pi/512
   cos[499]  =  15'b110000000011010;     //499pi/512
   sin[500]  =  15'b111110110100101;     //500pi/512
   cos[500]  =  15'b110000000010110;     //500pi/512
   sin[501]  =  15'b111110111010111;     //501pi/512
   cos[501]  =  15'b110000000010011;     //501pi/512
   sin[502]  =  15'b111111000001010;     //502pi/512
   cos[502]  =  15'b110000000001111;     //502pi/512
   sin[503]  =  15'b111111000111100;     //503pi/512
   cos[503]  =  15'b110000000001100;     //503pi/512
   sin[504]  =  15'b111111001101110;     //504pi/512
   cos[504]  =  15'b110000000001010;     //504pi/512
   sin[505]  =  15'b111111010100000;     //505pi/512
   cos[505]  =  15'b110000000001000;     //505pi/512
   sin[506]  =  15'b111111011010010;     //506pi/512
   cos[506]  =  15'b110000000000110;     //506pi/512
   sin[507]  =  15'b111111100000101;     //507pi/512
   cos[507]  =  15'b110000000000100;     //507pi/512
   sin[508]  =  15'b111111100110111;     //508pi/512
   cos[508]  =  15'b110000000000010;     //508pi/512
   sin[509]  =  15'b111111101101001;     //509pi/512
   cos[509]  =  15'b110000000000001;     //509pi/512
   sin[510]  =  15'b111111110011011;     //510pi/512
   cos[510]  =  15'b110000000000001;     //510pi/512
   sin[511]  =  15'b111111111001110;     //511pi/512
   cos[511]  =  15'b110000000000000;     //511pi/512
   m_sin[0]  =  15'b000000000000000;     //0pi/512
   m_cos[0]  =  15'b010000000000000;     //0pi/512
   m_sin[1]  =  15'b111111111011000;     //1pi/512
   m_cos[1]  =  15'b001111111111111;     //1pi/512
   m_sin[2]  =  15'b111111110110000;     //2pi/512
   m_cos[2]  =  15'b001111111111111;     //2pi/512
   m_sin[3]  =  15'b111111110000111;     //3pi/512
   m_cos[3]  =  15'b001111111111111;     //3pi/512
   m_sin[4]  =  15'b111111101011111;     //4pi/512
   m_cos[4]  =  15'b001111111111110;     //4pi/512
   m_sin[5]  =  15'b111111100110111;     //5pi/512
   m_cos[5]  =  15'b001111111111101;     //5pi/512
   m_sin[6]  =  15'b111111100001111;     //6pi/512
   m_cos[6]  =  15'b001111111111100;     //6pi/512
   m_sin[7]  =  15'b111111011100111;     //7pi/512
   m_cos[7]  =  15'b001111111111011;     //7pi/512
   m_sin[8]  =  15'b111111010111110;     //8pi/512
   m_cos[8]  =  15'b001111111111001;     //8pi/512
   m_sin[9]  =  15'b111111010010110;     //9pi/512
   m_cos[9]  =  15'b001111111111000;     //9pi/512
   m_sin[10]  =  15'b111111001101110;     //10pi/512
   m_cos[10]  =  15'b001111111110110;     //10pi/512
   m_sin[11]  =  15'b111111001000110;     //11pi/512
   m_cos[11]  =  15'b001111111110100;     //11pi/512
   m_sin[12]  =  15'b111111000011110;     //12pi/512
   m_cos[12]  =  15'b001111111110001;     //12pi/512
   m_sin[13]  =  15'b111110111110110;     //13pi/512
   m_cos[13]  =  15'b001111111101111;     //13pi/512
   m_sin[14]  =  15'b111110111001101;     //14pi/512
   m_cos[14]  =  15'b001111111101100;     //14pi/512
   m_sin[15]  =  15'b111110110100101;     //15pi/512
   m_cos[15]  =  15'b001111111101001;     //15pi/512
   m_sin[16]  =  15'b111110101111101;     //16pi/512
   m_cos[16]  =  15'b001111111100110;     //16pi/512
   m_sin[17]  =  15'b111110101010101;     //17pi/512
   m_cos[17]  =  15'b001111111100011;     //17pi/512
   m_sin[18]  =  15'b111110100101101;     //18pi/512
   m_cos[18]  =  15'b001111111100000;     //18pi/512
   m_sin[19]  =  15'b111110100000101;     //19pi/512
   m_cos[19]  =  15'b001111111011100;     //19pi/512
   m_sin[20]  =  15'b111110011011101;     //20pi/512
   m_cos[20]  =  15'b001111111011000;     //20pi/512
   m_sin[21]  =  15'b111110010110101;     //21pi/512
   m_cos[21]  =  15'b001111111010100;     //21pi/512
   m_sin[22]  =  15'b111110010001101;     //22pi/512
   m_cos[22]  =  15'b001111111010000;     //22pi/512
   m_sin[23]  =  15'b111110001100101;     //23pi/512
   m_cos[23]  =  15'b001111111001011;     //23pi/512
   m_sin[24]  =  15'b111110000111101;     //24pi/512
   m_cos[24]  =  15'b001111111000111;     //24pi/512
   m_sin[25]  =  15'b111110000010101;     //25pi/512
   m_cos[25]  =  15'b001111111000010;     //25pi/512
   m_sin[26]  =  15'b111101111101101;     //26pi/512
   m_cos[26]  =  15'b001111110111101;     //26pi/512
   m_sin[27]  =  15'b111101111000101;     //27pi/512
   m_cos[27]  =  15'b001111110111000;     //27pi/512
   m_sin[28]  =  15'b111101110011110;     //28pi/512
   m_cos[28]  =  15'b001111110110010;     //28pi/512
   m_sin[29]  =  15'b111101101110110;     //29pi/512
   m_cos[29]  =  15'b001111110101101;     //29pi/512
   m_sin[30]  =  15'b111101101001110;     //30pi/512
   m_cos[30]  =  15'b001111110100111;     //30pi/512
   m_sin[31]  =  15'b111101100100110;     //31pi/512
   m_cos[31]  =  15'b001111110100001;     //31pi/512
   m_sin[32]  =  15'b111101011111110;     //32pi/512
   m_cos[32]  =  15'b001111110011011;     //32pi/512
   m_sin[33]  =  15'b111101011010111;     //33pi/512
   m_cos[33]  =  15'b001111110010100;     //33pi/512
   m_sin[34]  =  15'b111101010101111;     //34pi/512
   m_cos[34]  =  15'b001111110001110;     //34pi/512
   m_sin[35]  =  15'b111101010000111;     //35pi/512
   m_cos[35]  =  15'b001111110000111;     //35pi/512
   m_sin[36]  =  15'b111101001100000;     //36pi/512
   m_cos[36]  =  15'b001111110000000;     //36pi/512
   m_sin[37]  =  15'b111101000111000;     //37pi/512
   m_cos[37]  =  15'b001111101111001;     //37pi/512
   m_sin[38]  =  15'b111101000010001;     //38pi/512
   m_cos[38]  =  15'b001111101110001;     //38pi/512
   m_sin[39]  =  15'b111100111101001;     //39pi/512
   m_cos[39]  =  15'b001111101101010;     //39pi/512
   m_sin[40]  =  15'b111100111000010;     //40pi/512
   m_cos[40]  =  15'b001111101100010;     //40pi/512
   m_sin[41]  =  15'b111100110011010;     //41pi/512
   m_cos[41]  =  15'b001111101011010;     //41pi/512
   m_sin[42]  =  15'b111100101110011;     //42pi/512
   m_cos[42]  =  15'b001111101010010;     //42pi/512
   m_sin[43]  =  15'b111100101001100;     //43pi/512
   m_cos[43]  =  15'b001111101001010;     //43pi/512
   m_sin[44]  =  15'b111100100100100;     //44pi/512
   m_cos[44]  =  15'b001111101000001;     //44pi/512
   m_sin[45]  =  15'b111100011111101;     //45pi/512
   m_cos[45]  =  15'b001111100111000;     //45pi/512
   m_sin[46]  =  15'b111100011010110;     //46pi/512
   m_cos[46]  =  15'b001111100110000;     //46pi/512
   m_sin[47]  =  15'b111100010101111;     //47pi/512
   m_cos[47]  =  15'b001111100100110;     //47pi/512
   m_sin[48]  =  15'b111100010001000;     //48pi/512
   m_cos[48]  =  15'b001111100011101;     //48pi/512
   m_sin[49]  =  15'b111100001100001;     //49pi/512
   m_cos[49]  =  15'b001111100010100;     //49pi/512
   m_sin[50]  =  15'b111100000111010;     //50pi/512
   m_cos[50]  =  15'b001111100001010;     //50pi/512
   m_sin[51]  =  15'b111100000010011;     //51pi/512
   m_cos[51]  =  15'b001111100000000;     //51pi/512
   m_sin[52]  =  15'b111011111101100;     //52pi/512
   m_cos[52]  =  15'b001111011110110;     //52pi/512
   m_sin[53]  =  15'b111011111000101;     //53pi/512
   m_cos[53]  =  15'b001111011101100;     //53pi/512
   m_sin[54]  =  15'b111011110011110;     //54pi/512
   m_cos[54]  =  15'b001111011100001;     //54pi/512
   m_sin[55]  =  15'b111011101110111;     //55pi/512
   m_cos[55]  =  15'b001111011010111;     //55pi/512
   m_sin[56]  =  15'b111011101010000;     //56pi/512
   m_cos[56]  =  15'b001111011001100;     //56pi/512
   m_sin[57]  =  15'b111011100101010;     //57pi/512
   m_cos[57]  =  15'b001111011000001;     //57pi/512
   m_sin[58]  =  15'b111011100000011;     //58pi/512
   m_cos[58]  =  15'b001111010110110;     //58pi/512
   m_sin[59]  =  15'b111011011011100;     //59pi/512
   m_cos[59]  =  15'b001111010101010;     //59pi/512
   m_sin[60]  =  15'b111011010110110;     //60pi/512
   m_cos[60]  =  15'b001111010011111;     //60pi/512
   m_sin[61]  =  15'b111011010010000;     //61pi/512
   m_cos[61]  =  15'b001111010010011;     //61pi/512
   m_sin[62]  =  15'b111011001101001;     //62pi/512
   m_cos[62]  =  15'b001111010000111;     //62pi/512
   m_sin[63]  =  15'b111011001000011;     //63pi/512
   m_cos[63]  =  15'b001111001111011;     //63pi/512
   m_sin[64]  =  15'b111011000011101;     //64pi/512
   m_cos[64]  =  15'b001111001101111;     //64pi/512
   m_sin[65]  =  15'b111010111110110;     //65pi/512
   m_cos[65]  =  15'b001111001100010;     //65pi/512
   m_sin[66]  =  15'b111010111010000;     //66pi/512
   m_cos[66]  =  15'b001111001010101;     //66pi/512
   m_sin[67]  =  15'b111010110101010;     //67pi/512
   m_cos[67]  =  15'b001111001001000;     //67pi/512
   m_sin[68]  =  15'b111010110000100;     //68pi/512
   m_cos[68]  =  15'b001111000111011;     //68pi/512
   m_sin[69]  =  15'b111010101011110;     //69pi/512
   m_cos[69]  =  15'b001111000101110;     //69pi/512
   m_sin[70]  =  15'b111010100111000;     //70pi/512
   m_cos[70]  =  15'b001111000100001;     //70pi/512
   m_sin[71]  =  15'b111010100010010;     //71pi/512
   m_cos[71]  =  15'b001111000010011;     //71pi/512
   m_sin[72]  =  15'b111010011101101;     //72pi/512
   m_cos[72]  =  15'b001111000000101;     //72pi/512
   m_sin[73]  =  15'b111010011000111;     //73pi/512
   m_cos[73]  =  15'b001110111110111;     //73pi/512
   m_sin[74]  =  15'b111010010100001;     //74pi/512
   m_cos[74]  =  15'b001110111101001;     //74pi/512
   m_sin[75]  =  15'b111010001111100;     //75pi/512
   m_cos[75]  =  15'b001110111011011;     //75pi/512
   m_sin[76]  =  15'b111010001010110;     //76pi/512
   m_cos[76]  =  15'b001110111001100;     //76pi/512
   m_sin[77]  =  15'b111010000110001;     //77pi/512
   m_cos[77]  =  15'b001110110111101;     //77pi/512
   m_sin[78]  =  15'b111010000001100;     //78pi/512
   m_cos[78]  =  15'b001110110101110;     //78pi/512
   m_sin[79]  =  15'b111001111100110;     //79pi/512
   m_cos[79]  =  15'b001110110011111;     //79pi/512
   m_sin[80]  =  15'b111001111000001;     //80pi/512
   m_cos[80]  =  15'b001110110010000;     //80pi/512
   m_sin[81]  =  15'b111001110011100;     //81pi/512
   m_cos[81]  =  15'b001110110000000;     //81pi/512
   m_sin[82]  =  15'b111001101110111;     //82pi/512
   m_cos[82]  =  15'b001110101110001;     //82pi/512
   m_sin[83]  =  15'b111001101010010;     //83pi/512
   m_cos[83]  =  15'b001110101100001;     //83pi/512
   m_sin[84]  =  15'b111001100101101;     //84pi/512
   m_cos[84]  =  15'b001110101010001;     //84pi/512
   m_sin[85]  =  15'b111001100001000;     //85pi/512
   m_cos[85]  =  15'b001110101000001;     //85pi/512
   m_sin[86]  =  15'b111001011100100;     //86pi/512
   m_cos[86]  =  15'b001110100110000;     //86pi/512
   m_sin[87]  =  15'b111001010111111;     //87pi/512
   m_cos[87]  =  15'b001110100100000;     //87pi/512
   m_sin[88]  =  15'b111001010011010;     //88pi/512
   m_cos[88]  =  15'b001110100001111;     //88pi/512
   m_sin[89]  =  15'b111001001110110;     //89pi/512
   m_cos[89]  =  15'b001110011111110;     //89pi/512
   m_sin[90]  =  15'b111001001010001;     //90pi/512
   m_cos[90]  =  15'b001110011101101;     //90pi/512
   m_sin[91]  =  15'b111001000101101;     //91pi/512
   m_cos[91]  =  15'b001110011011100;     //91pi/512
   m_sin[92]  =  15'b111001000001001;     //92pi/512
   m_cos[92]  =  15'b001110011001010;     //92pi/512
   m_sin[93]  =  15'b111000111100101;     //93pi/512
   m_cos[93]  =  15'b001110010111001;     //93pi/512
   m_sin[94]  =  15'b111000111000001;     //94pi/512
   m_cos[94]  =  15'b001110010100111;     //94pi/512
   m_sin[95]  =  15'b111000110011101;     //95pi/512
   m_cos[95]  =  15'b001110010010101;     //95pi/512
   m_sin[96]  =  15'b111000101111001;     //96pi/512
   m_cos[96]  =  15'b001110010000011;     //96pi/512
   m_sin[97]  =  15'b111000101010101;     //97pi/512
   m_cos[97]  =  15'b001110001110000;     //97pi/512
   m_sin[98]  =  15'b111000100110001;     //98pi/512
   m_cos[98]  =  15'b001110001011110;     //98pi/512
   m_sin[99]  =  15'b111000100001110;     //99pi/512
   m_cos[99]  =  15'b001110001001011;     //99pi/512
   m_sin[100]  =  15'b111000011101010;     //100pi/512
   m_cos[100]  =  15'b001110000111000;     //100pi/512
   m_sin[101]  =  15'b111000011000111;     //101pi/512
   m_cos[101]  =  15'b001110000100101;     //101pi/512
   m_sin[102]  =  15'b111000010100100;     //102pi/512
   m_cos[102]  =  15'b001110000010010;     //102pi/512
   m_sin[103]  =  15'b111000010000000;     //103pi/512
   m_cos[103]  =  15'b001101111111111;     //103pi/512
   m_sin[104]  =  15'b111000001011101;     //104pi/512
   m_cos[104]  =  15'b001101111101011;     //104pi/512
   m_sin[105]  =  15'b111000000111010;     //105pi/512
   m_cos[105]  =  15'b001101111010111;     //105pi/512
   m_sin[106]  =  15'b111000000010111;     //106pi/512
   m_cos[106]  =  15'b001101111000011;     //106pi/512
   m_sin[107]  =  15'b110111111110100;     //107pi/512
   m_cos[107]  =  15'b001101110101111;     //107pi/512
   m_sin[108]  =  15'b110111111010010;     //108pi/512
   m_cos[108]  =  15'b001101110011011;     //108pi/512
   m_sin[109]  =  15'b110111110101111;     //109pi/512
   m_cos[109]  =  15'b001101110000111;     //109pi/512
   m_sin[110]  =  15'b110111110001100;     //110pi/512
   m_cos[110]  =  15'b001101101110010;     //110pi/512
   m_sin[111]  =  15'b110111101101010;     //111pi/512
   m_cos[111]  =  15'b001101101011101;     //111pi/512
   m_sin[112]  =  15'b110111101001000;     //112pi/512
   m_cos[112]  =  15'b001101101001000;     //112pi/512
   m_sin[113]  =  15'b110111100100101;     //113pi/512
   m_cos[113]  =  15'b001101100110011;     //113pi/512
   m_sin[114]  =  15'b110111100000011;     //114pi/512
   m_cos[114]  =  15'b001101100011110;     //114pi/512
   m_sin[115]  =  15'b110111011100001;     //115pi/512
   m_cos[115]  =  15'b001101100001001;     //115pi/512
   m_sin[116]  =  15'b110111010111111;     //116pi/512
   m_cos[116]  =  15'b001101011110011;     //116pi/512
   m_sin[117]  =  15'b110111010011110;     //117pi/512
   m_cos[117]  =  15'b001101011011101;     //117pi/512
   m_sin[118]  =  15'b110111001111100;     //118pi/512
   m_cos[118]  =  15'b001101011000111;     //118pi/512
   m_sin[119]  =  15'b110111001011010;     //119pi/512
   m_cos[119]  =  15'b001101010110001;     //119pi/512
   m_sin[120]  =  15'b110111000111001;     //120pi/512
   m_cos[120]  =  15'b001101010011011;     //120pi/512
   m_sin[121]  =  15'b110111000010111;     //121pi/512
   m_cos[121]  =  15'b001101010000100;     //121pi/512
   m_sin[122]  =  15'b110110111110110;     //122pi/512
   m_cos[122]  =  15'b001101001101110;     //122pi/512
   m_sin[123]  =  15'b110110111010101;     //123pi/512
   m_cos[123]  =  15'b001101001010111;     //123pi/512
   m_sin[124]  =  15'b110110110110100;     //124pi/512
   m_cos[124]  =  15'b001101001000000;     //124pi/512
   m_sin[125]  =  15'b110110110010011;     //125pi/512
   m_cos[125]  =  15'b001101000101001;     //125pi/512
   m_sin[126]  =  15'b110110101110010;     //126pi/512
   m_cos[126]  =  15'b001101000010010;     //126pi/512
   m_sin[127]  =  15'b110110101010001;     //127pi/512
   m_cos[127]  =  15'b001100111111011;     //127pi/512
   m_sin[128]  =  15'b110110100110001;     //128pi/512
   m_cos[128]  =  15'b001100111100011;     //128pi/512
   m_sin[129]  =  15'b110110100010000;     //129pi/512
   m_cos[129]  =  15'b001100111001011;     //129pi/512
   m_sin[130]  =  15'b110110011110000;     //130pi/512
   m_cos[130]  =  15'b001100110110011;     //130pi/512
   m_sin[131]  =  15'b110110011010000;     //131pi/512
   m_cos[131]  =  15'b001100110011011;     //131pi/512
   m_sin[132]  =  15'b110110010110000;     //132pi/512
   m_cos[132]  =  15'b001100110000011;     //132pi/512
   m_sin[133]  =  15'b110110010010000;     //133pi/512
   m_cos[133]  =  15'b001100101101011;     //133pi/512
   m_sin[134]  =  15'b110110001110000;     //134pi/512
   m_cos[134]  =  15'b001100101010010;     //134pi/512
   m_sin[135]  =  15'b110110001010000;     //135pi/512
   m_cos[135]  =  15'b001100100111010;     //135pi/512
   m_sin[136]  =  15'b110110000110000;     //136pi/512
   m_cos[136]  =  15'b001100100100001;     //136pi/512
   m_sin[137]  =  15'b110110000010001;     //137pi/512
   m_cos[137]  =  15'b001100100001000;     //137pi/512
   m_sin[138]  =  15'b110101111110001;     //138pi/512
   m_cos[138]  =  15'b001100011101111;     //138pi/512
   m_sin[139]  =  15'b110101111010010;     //139pi/512
   m_cos[139]  =  15'b001100011010101;     //139pi/512
   m_sin[140]  =  15'b110101110110011;     //140pi/512
   m_cos[140]  =  15'b001100010111100;     //140pi/512
   m_sin[141]  =  15'b110101110010100;     //141pi/512
   m_cos[141]  =  15'b001100010100010;     //141pi/512
   m_sin[142]  =  15'b110101101110101;     //142pi/512
   m_cos[142]  =  15'b001100010001001;     //142pi/512
   m_sin[143]  =  15'b110101101010110;     //143pi/512
   m_cos[143]  =  15'b001100001101111;     //143pi/512
   m_sin[144]  =  15'b110101100111000;     //144pi/512
   m_cos[144]  =  15'b001100001010101;     //144pi/512
   m_sin[145]  =  15'b110101100011001;     //145pi/512
   m_cos[145]  =  15'b001100000111011;     //145pi/512
   m_sin[146]  =  15'b110101011111011;     //146pi/512
   m_cos[146]  =  15'b001100000100000;     //146pi/512
   m_sin[147]  =  15'b110101011011101;     //147pi/512
   m_cos[147]  =  15'b001100000000110;     //147pi/512
   m_sin[148]  =  15'b110101010111110;     //148pi/512
   m_cos[148]  =  15'b001011111101011;     //148pi/512
   m_sin[149]  =  15'b110101010100000;     //149pi/512
   m_cos[149]  =  15'b001011111010000;     //149pi/512
   m_sin[150]  =  15'b110101010000011;     //150pi/512
   m_cos[150]  =  15'b001011110110101;     //150pi/512
   m_sin[151]  =  15'b110101001100101;     //151pi/512
   m_cos[151]  =  15'b001011110011010;     //151pi/512
   m_sin[152]  =  15'b110101001000111;     //152pi/512
   m_cos[152]  =  15'b001011101111111;     //152pi/512
   m_sin[153]  =  15'b110101000101010;     //153pi/512
   m_cos[153]  =  15'b001011101100100;     //153pi/512
   m_sin[154]  =  15'b110101000001100;     //154pi/512
   m_cos[154]  =  15'b001011101001000;     //154pi/512
   m_sin[155]  =  15'b110100111101111;     //155pi/512
   m_cos[155]  =  15'b001011100101101;     //155pi/512
   m_sin[156]  =  15'b110100111010010;     //156pi/512
   m_cos[156]  =  15'b001011100010001;     //156pi/512
   m_sin[157]  =  15'b110100110110101;     //157pi/512
   m_cos[157]  =  15'b001011011110101;     //157pi/512
   m_sin[158]  =  15'b110100110011001;     //158pi/512
   m_cos[158]  =  15'b001011011011001;     //158pi/512
   m_sin[159]  =  15'b110100101111100;     //159pi/512
   m_cos[159]  =  15'b001011010111100;     //159pi/512
   m_sin[160]  =  15'b110100101011111;     //160pi/512
   m_cos[160]  =  15'b001011010100000;     //160pi/512
   m_sin[161]  =  15'b110100101000011;     //161pi/512
   m_cos[161]  =  15'b001011010000100;     //161pi/512
   m_sin[162]  =  15'b110100100100111;     //162pi/512
   m_cos[162]  =  15'b001011001100111;     //162pi/512
   m_sin[163]  =  15'b110100100001011;     //163pi/512
   m_cos[163]  =  15'b001011001001010;     //163pi/512
   m_sin[164]  =  15'b110100011101111;     //164pi/512
   m_cos[164]  =  15'b001011000101101;     //164pi/512
   m_sin[165]  =  15'b110100011010011;     //165pi/512
   m_cos[165]  =  15'b001011000010000;     //165pi/512
   m_sin[166]  =  15'b110100010110111;     //166pi/512
   m_cos[166]  =  15'b001010111110011;     //166pi/512
   m_sin[167]  =  15'b110100010011100;     //167pi/512
   m_cos[167]  =  15'b001010111010110;     //167pi/512
   m_sin[168]  =  15'b110100010000000;     //168pi/512
   m_cos[168]  =  15'b001010110111000;     //168pi/512
   m_sin[169]  =  15'b110100001100101;     //169pi/512
   m_cos[169]  =  15'b001010110011011;     //169pi/512
   m_sin[170]  =  15'b110100001001010;     //170pi/512
   m_cos[170]  =  15'b001010101111101;     //170pi/512
   m_sin[171]  =  15'b110100000101111;     //171pi/512
   m_cos[171]  =  15'b001010101011111;     //171pi/512
   m_sin[172]  =  15'b110100000010100;     //172pi/512
   m_cos[172]  =  15'b001010101000001;     //172pi/512
   m_sin[173]  =  15'b110011111111010;     //173pi/512
   m_cos[173]  =  15'b001010100100011;     //173pi/512
   m_sin[174]  =  15'b110011111011111;     //174pi/512
   m_cos[174]  =  15'b001010100000101;     //174pi/512
   m_sin[175]  =  15'b110011111000101;     //175pi/512
   m_cos[175]  =  15'b001010011100110;     //175pi/512
   m_sin[176]  =  15'b110011110101011;     //176pi/512
   m_cos[176]  =  15'b001010011001000;     //176pi/512
   m_sin[177]  =  15'b110011110010001;     //177pi/512
   m_cos[177]  =  15'b001010010101001;     //177pi/512
   m_sin[178]  =  15'b110011101110111;     //178pi/512
   m_cos[178]  =  15'b001010010001010;     //178pi/512
   m_sin[179]  =  15'b110011101011101;     //179pi/512
   m_cos[179]  =  15'b001010001101011;     //179pi/512
   m_sin[180]  =  15'b110011101000011;     //180pi/512
   m_cos[180]  =  15'b001010001001100;     //180pi/512
   m_sin[181]  =  15'b110011100101010;     //181pi/512
   m_cos[181]  =  15'b001010000101101;     //181pi/512
   m_sin[182]  =  15'b110011100010001;     //182pi/512
   m_cos[182]  =  15'b001010000001110;     //182pi/512
   m_sin[183]  =  15'b110011011111000;     //183pi/512
   m_cos[183]  =  15'b001001111101111;     //183pi/512
   m_sin[184]  =  15'b110011011011111;     //184pi/512
   m_cos[184]  =  15'b001001111001111;     //184pi/512
   m_sin[185]  =  15'b110011011000110;     //185pi/512
   m_cos[185]  =  15'b001001110101111;     //185pi/512
   m_sin[186]  =  15'b110011010101101;     //186pi/512
   m_cos[186]  =  15'b001001110010000;     //186pi/512
   m_sin[187]  =  15'b110011010010101;     //187pi/512
   m_cos[187]  =  15'b001001101110000;     //187pi/512
   m_sin[188]  =  15'b110011001111100;     //188pi/512
   m_cos[188]  =  15'b001001101010000;     //188pi/512
   m_sin[189]  =  15'b110011001100100;     //189pi/512
   m_cos[189]  =  15'b001001100110000;     //189pi/512
   m_sin[190]  =  15'b110011001001100;     //190pi/512
   m_cos[190]  =  15'b001001100001111;     //190pi/512
   m_sin[191]  =  15'b110011000110100;     //191pi/512
   m_cos[191]  =  15'b001001011101111;     //191pi/512
   m_sin[192]  =  15'b110011000011101;     //192pi/512
   m_cos[192]  =  15'b001001011001111;     //192pi/512
   m_sin[193]  =  15'b110011000000101;     //193pi/512
   m_cos[193]  =  15'b001001010101110;     //193pi/512
   m_sin[194]  =  15'b110010111101110;     //194pi/512
   m_cos[194]  =  15'b001001010001101;     //194pi/512
   m_sin[195]  =  15'b110010111010110;     //195pi/512
   m_cos[195]  =  15'b001001001101101;     //195pi/512
   m_sin[196]  =  15'b110010110111111;     //196pi/512
   m_cos[196]  =  15'b001001001001100;     //196pi/512
   m_sin[197]  =  15'b110010110101000;     //197pi/512
   m_cos[197]  =  15'b001001000101011;     //197pi/512
   m_sin[198]  =  15'b110010110010010;     //198pi/512
   m_cos[198]  =  15'b001001000001001;     //198pi/512
   m_sin[199]  =  15'b110010101111011;     //199pi/512
   m_cos[199]  =  15'b001000111101000;     //199pi/512
   m_sin[200]  =  15'b110010101100101;     //200pi/512
   m_cos[200]  =  15'b001000111000111;     //200pi/512
   m_sin[201]  =  15'b110010101001110;     //201pi/512
   m_cos[201]  =  15'b001000110100101;     //201pi/512
   m_sin[202]  =  15'b110010100111000;     //202pi/512
   m_cos[202]  =  15'b001000110000100;     //202pi/512
   m_sin[203]  =  15'b110010100100010;     //203pi/512
   m_cos[203]  =  15'b001000101100010;     //203pi/512
   m_sin[204]  =  15'b110010100001101;     //204pi/512
   m_cos[204]  =  15'b001000101000000;     //204pi/512
   m_sin[205]  =  15'b110010011110111;     //205pi/512
   m_cos[205]  =  15'b001000100011110;     //205pi/512
   m_sin[206]  =  15'b110010011100010;     //206pi/512
   m_cos[206]  =  15'b001000011111100;     //206pi/512
   m_sin[207]  =  15'b110010011001100;     //207pi/512
   m_cos[207]  =  15'b001000011011010;     //207pi/512
   m_sin[208]  =  15'b110010010110111;     //208pi/512
   m_cos[208]  =  15'b001000010111000;     //208pi/512
   m_sin[209]  =  15'b110010010100010;     //209pi/512
   m_cos[209]  =  15'b001000010010101;     //209pi/512
   m_sin[210]  =  15'b110010010001101;     //210pi/512
   m_cos[210]  =  15'b001000001110011;     //210pi/512
   m_sin[211]  =  15'b110010001111001;     //211pi/512
   m_cos[211]  =  15'b001000001010000;     //211pi/512
   m_sin[212]  =  15'b110010001100100;     //212pi/512
   m_cos[212]  =  15'b001000000101110;     //212pi/512
   m_sin[213]  =  15'b110010001010000;     //213pi/512
   m_cos[213]  =  15'b001000000001011;     //213pi/512
   m_sin[214]  =  15'b110010000111100;     //214pi/512
   m_cos[214]  =  15'b000111111101000;     //214pi/512
   m_sin[215]  =  15'b110010000101000;     //215pi/512
   m_cos[215]  =  15'b000111111000101;     //215pi/512
   m_sin[216]  =  15'b110010000010101;     //216pi/512
   m_cos[216]  =  15'b000111110100010;     //216pi/512
   m_sin[217]  =  15'b110010000000001;     //217pi/512
   m_cos[217]  =  15'b000111101111111;     //217pi/512
   m_sin[218]  =  15'b110001111101110;     //218pi/512
   m_cos[218]  =  15'b000111101011100;     //218pi/512
   m_sin[219]  =  15'b110001111011010;     //219pi/512
   m_cos[219]  =  15'b000111100111001;     //219pi/512
   m_sin[220]  =  15'b110001111000111;     //220pi/512
   m_cos[220]  =  15'b000111100010101;     //220pi/512
   m_sin[221]  =  15'b110001110110100;     //221pi/512
   m_cos[221]  =  15'b000111011110010;     //221pi/512
   m_sin[222]  =  15'b110001110100010;     //222pi/512
   m_cos[222]  =  15'b000111011001110;     //222pi/512
   m_sin[223]  =  15'b110001110001111;     //223pi/512
   m_cos[223]  =  15'b000111010101010;     //223pi/512
   m_sin[224]  =  15'b110001101111101;     //224pi/512
   m_cos[224]  =  15'b000111010000111;     //224pi/512
   m_sin[225]  =  15'b110001101101011;     //225pi/512
   m_cos[225]  =  15'b000111001100011;     //225pi/512
   m_sin[226]  =  15'b110001101011001;     //226pi/512
   m_cos[226]  =  15'b000111000111111;     //226pi/512
   m_sin[227]  =  15'b110001101000111;     //227pi/512
   m_cos[227]  =  15'b000111000011011;     //227pi/512
   m_sin[228]  =  15'b110001100110101;     //228pi/512
   m_cos[228]  =  15'b000110111110111;     //228pi/512
   m_sin[229]  =  15'b110001100100100;     //229pi/512
   m_cos[229]  =  15'b000110111010010;     //229pi/512
   m_sin[230]  =  15'b110001100010011;     //230pi/512
   m_cos[230]  =  15'b000110110101110;     //230pi/512
   m_sin[231]  =  15'b110001100000001;     //231pi/512
   m_cos[231]  =  15'b000110110001010;     //231pi/512
   m_sin[232]  =  15'b110001011110000;     //232pi/512
   m_cos[232]  =  15'b000110101100101;     //232pi/512
   m_sin[233]  =  15'b110001011100000;     //233pi/512
   m_cos[233]  =  15'b000110101000001;     //233pi/512
   m_sin[234]  =  15'b110001011001111;     //234pi/512
   m_cos[234]  =  15'b000110100011100;     //234pi/512
   m_sin[235]  =  15'b110001010111111;     //235pi/512
   m_cos[235]  =  15'b000110011110111;     //235pi/512
   m_sin[236]  =  15'b110001010101111;     //236pi/512
   m_cos[236]  =  15'b000110011010010;     //236pi/512
   m_sin[237]  =  15'b110001010011111;     //237pi/512
   m_cos[237]  =  15'b000110010101110;     //237pi/512
   m_sin[238]  =  15'b110001010001111;     //238pi/512
   m_cos[238]  =  15'b000110010001001;     //238pi/512
   m_sin[239]  =  15'b110001001111111;     //239pi/512
   m_cos[239]  =  15'b000110001100100;     //239pi/512
   m_sin[240]  =  15'b110001001110000;     //240pi/512
   m_cos[240]  =  15'b000110000111110;     //240pi/512
   m_sin[241]  =  15'b110001001100000;     //241pi/512
   m_cos[241]  =  15'b000110000011001;     //241pi/512
   m_sin[242]  =  15'b110001001010001;     //242pi/512
   m_cos[242]  =  15'b000101111110100;     //242pi/512
   m_sin[243]  =  15'b110001001000010;     //243pi/512
   m_cos[243]  =  15'b000101111001111;     //243pi/512
   m_sin[244]  =  15'b110001000110011;     //244pi/512
   m_cos[244]  =  15'b000101110101001;     //244pi/512
   m_sin[245]  =  15'b110001000100101;     //245pi/512
   m_cos[245]  =  15'b000101110000100;     //245pi/512
   m_sin[246]  =  15'b110001000010111;     //246pi/512
   m_cos[246]  =  15'b000101101011110;     //246pi/512
   m_sin[247]  =  15'b110001000001000;     //247pi/512
   m_cos[247]  =  15'b000101100111001;     //247pi/512
   m_sin[248]  =  15'b110000111111010;     //248pi/512
   m_cos[248]  =  15'b000101100010011;     //248pi/512
   m_sin[249]  =  15'b110000111101101;     //249pi/512
   m_cos[249]  =  15'b000101011101101;     //249pi/512
   m_sin[250]  =  15'b110000111011111;     //250pi/512
   m_cos[250]  =  15'b000101011000111;     //250pi/512
   m_sin[251]  =  15'b110000111010001;     //251pi/512
   m_cos[251]  =  15'b000101010100001;     //251pi/512
   m_sin[252]  =  15'b110000111000100;     //252pi/512
   m_cos[252]  =  15'b000101001111011;     //252pi/512
   m_sin[253]  =  15'b110000110110111;     //253pi/512
   m_cos[253]  =  15'b000101001010101;     //253pi/512
   m_sin[254]  =  15'b110000110101010;     //254pi/512
   m_cos[254]  =  15'b000101000101111;     //254pi/512
   m_sin[255]  =  15'b110000110011101;     //255pi/512
   m_cos[255]  =  15'b000101000001001;     //255pi/512
   m_sin[256]  =  15'b110000110010001;     //256pi/512
   m_cos[256]  =  15'b000100111100011;     //256pi/512
   m_sin[257]  =  15'b110000110000101;     //257pi/512
   m_cos[257]  =  15'b000100110111101;     //257pi/512
   m_sin[258]  =  15'b110000101111000;     //258pi/512
   m_cos[258]  =  15'b000100110010110;     //258pi/512
   m_sin[259]  =  15'b110000101101101;     //259pi/512
   m_cos[259]  =  15'b000100101110000;     //259pi/512
   m_sin[260]  =  15'b110000101100001;     //260pi/512
   m_cos[260]  =  15'b000100101001010;     //260pi/512
   m_sin[261]  =  15'b110000101010101;     //261pi/512
   m_cos[261]  =  15'b000100100100011;     //261pi/512
   m_sin[262]  =  15'b110000101001010;     //262pi/512
   m_cos[262]  =  15'b000100011111100;     //262pi/512
   m_sin[263]  =  15'b110000100111111;     //263pi/512
   m_cos[263]  =  15'b000100011010110;     //263pi/512
   m_sin[264]  =  15'b110000100110100;     //264pi/512
   m_cos[264]  =  15'b000100010101111;     //264pi/512
   m_sin[265]  =  15'b110000100101001;     //265pi/512
   m_cos[265]  =  15'b000100010001000;     //265pi/512
   m_sin[266]  =  15'b110000100011110;     //266pi/512
   m_cos[266]  =  15'b000100001100010;     //266pi/512
   m_sin[267]  =  15'b110000100010100;     //267pi/512
   m_cos[267]  =  15'b000100000111011;     //267pi/512
   m_sin[268]  =  15'b110000100001001;     //268pi/512
   m_cos[268]  =  15'b000100000010100;     //268pi/512
   m_sin[269]  =  15'b110000011111111;     //269pi/512
   m_cos[269]  =  15'b000011111101101;     //269pi/512
   m_sin[270]  =  15'b110000011110110;     //270pi/512
   m_cos[270]  =  15'b000011111000110;     //270pi/512
   m_sin[271]  =  15'b110000011101100;     //271pi/512
   m_cos[271]  =  15'b000011110011111;     //271pi/512
   m_sin[272]  =  15'b110000011100010;     //272pi/512
   m_cos[272]  =  15'b000011101111000;     //272pi/512
   m_sin[273]  =  15'b110000011011001;     //273pi/512
   m_cos[273]  =  15'b000011101010001;     //273pi/512
   m_sin[274]  =  15'b110000011010000;     //274pi/512
   m_cos[274]  =  15'b000011100101010;     //274pi/512
   m_sin[275]  =  15'b110000011000111;     //275pi/512
   m_cos[275]  =  15'b000011100000010;     //275pi/512
   m_sin[276]  =  15'b110000010111110;     //276pi/512
   m_cos[276]  =  15'b000011011011011;     //276pi/512
   m_sin[277]  =  15'b110000010110110;     //277pi/512
   m_cos[277]  =  15'b000011010110100;     //277pi/512
   m_sin[278]  =  15'b110000010101101;     //278pi/512
   m_cos[278]  =  15'b000011010001100;     //278pi/512
   m_sin[279]  =  15'b110000010100101;     //279pi/512
   m_cos[279]  =  15'b000011001100101;     //279pi/512
   m_sin[280]  =  15'b110000010011101;     //280pi/512
   m_cos[280]  =  15'b000011000111110;     //280pi/512
   m_sin[281]  =  15'b110000010010110;     //281pi/512
   m_cos[281]  =  15'b000011000010110;     //281pi/512
   m_sin[282]  =  15'b110000010001110;     //282pi/512
   m_cos[282]  =  15'b000010111101111;     //282pi/512
   m_sin[283]  =  15'b110000010000111;     //283pi/512
   m_cos[283]  =  15'b000010111000111;     //283pi/512
   m_sin[284]  =  15'b110000010000000;     //284pi/512
   m_cos[284]  =  15'b000010110100000;     //284pi/512
   m_sin[285]  =  15'b110000001111001;     //285pi/512
   m_cos[285]  =  15'b000010101111000;     //285pi/512
   m_sin[286]  =  15'b110000001110010;     //286pi/512
   m_cos[286]  =  15'b000010101010000;     //286pi/512
   m_sin[287]  =  15'b110000001101011;     //287pi/512
   m_cos[287]  =  15'b000010100101001;     //287pi/512
   m_sin[288]  =  15'b110000001100101;     //288pi/512
   m_cos[288]  =  15'b000010100000001;     //288pi/512
   m_sin[289]  =  15'b110000001011111;     //289pi/512
   m_cos[289]  =  15'b000010011011001;     //289pi/512
   m_sin[290]  =  15'b110000001011001;     //290pi/512
   m_cos[290]  =  15'b000010010110010;     //290pi/512
   m_sin[291]  =  15'b110000001010011;     //291pi/512
   m_cos[291]  =  15'b000010010001010;     //291pi/512
   m_sin[292]  =  15'b110000001001101;     //292pi/512
   m_cos[292]  =  15'b000010001100010;     //292pi/512
   m_sin[293]  =  15'b110000001001000;     //293pi/512
   m_cos[293]  =  15'b000010000111010;     //293pi/512
   m_sin[294]  =  15'b110000001000011;     //294pi/512
   m_cos[294]  =  15'b000010000010010;     //294pi/512
   m_sin[295]  =  15'b110000000111110;     //295pi/512
   m_cos[295]  =  15'b000001111101010;     //295pi/512
   m_sin[296]  =  15'b110000000111001;     //296pi/512
   m_cos[296]  =  15'b000001111000010;     //296pi/512
   m_sin[297]  =  15'b110000000110100;     //297pi/512
   m_cos[297]  =  15'b000001110011010;     //297pi/512
   m_sin[298]  =  15'b110000000110000;     //298pi/512
   m_cos[298]  =  15'b000001101110010;     //298pi/512
   m_sin[299]  =  15'b110000000101011;     //299pi/512
   m_cos[299]  =  15'b000001101001010;     //299pi/512
   m_sin[300]  =  15'b110000000100111;     //300pi/512
   m_cos[300]  =  15'b000001100100010;     //300pi/512
   m_sin[301]  =  15'b110000000100100;     //301pi/512
   m_cos[301]  =  15'b000001011111010;     //301pi/512
   m_sin[302]  =  15'b110000000100000;     //302pi/512
   m_cos[302]  =  15'b000001011010010;     //302pi/512
   m_sin[303]  =  15'b110000000011101;     //303pi/512
   m_cos[303]  =  15'b000001010101010;     //303pi/512
   m_sin[304]  =  15'b110000000011001;     //304pi/512
   m_cos[304]  =  15'b000001010000010;     //304pi/512
   m_sin[305]  =  15'b110000000010110;     //305pi/512
   m_cos[305]  =  15'b000001001011010;     //305pi/512
   m_sin[306]  =  15'b110000000010011;     //306pi/512
   m_cos[306]  =  15'b000001000110010;     //306pi/512
   m_sin[307]  =  15'b110000000010001;     //307pi/512
   m_cos[307]  =  15'b000001000001010;     //307pi/512
   m_sin[308]  =  15'b110000000001110;     //308pi/512
   m_cos[308]  =  15'b000000111100010;     //308pi/512
   m_sin[309]  =  15'b110000000001100;     //309pi/512
   m_cos[309]  =  15'b000000110111010;     //309pi/512
   m_sin[310]  =  15'b110000000001010;     //310pi/512
   m_cos[310]  =  15'b000000110010001;     //310pi/512
   m_sin[311]  =  15'b110000000001000;     //311pi/512
   m_cos[311]  =  15'b000000101101001;     //311pi/512
   m_sin[312]  =  15'b110000000000110;     //312pi/512
   m_cos[312]  =  15'b000000101000001;     //312pi/512
   m_sin[313]  =  15'b110000000000101;     //313pi/512
   m_cos[313]  =  15'b000000100011001;     //313pi/512
   m_sin[314]  =  15'b110000000000100;     //314pi/512
   m_cos[314]  =  15'b000000011110001;     //314pi/512
   m_sin[315]  =  15'b110000000000010;     //315pi/512
   m_cos[315]  =  15'b000000011001001;     //315pi/512
   m_sin[316]  =  15'b110000000000010;     //316pi/512
   m_cos[316]  =  15'b000000010100000;     //316pi/512
   m_sin[317]  =  15'b110000000000001;     //317pi/512
   m_cos[317]  =  15'b000000001111000;     //317pi/512
   m_sin[318]  =  15'b110000000000000;     //318pi/512
   m_cos[318]  =  15'b000000001010000;     //318pi/512
   m_sin[319]  =  15'b110000000000000;     //319pi/512
   m_cos[319]  =  15'b000000000101000;     //319pi/512
   m_sin[320]  =  15'b110000000000000;     //320pi/512
   m_cos[320]  =  15'b000000000000000;     //320pi/512
   m_sin[321]  =  15'b110000000000000;     //321pi/512
   m_cos[321]  =  15'b111111111011000;     //321pi/512
   m_sin[322]  =  15'b110000000000000;     //322pi/512
   m_cos[322]  =  15'b111111110110000;     //322pi/512
   m_sin[323]  =  15'b110000000000001;     //323pi/512
   m_cos[323]  =  15'b111111110000111;     //323pi/512
   m_sin[324]  =  15'b110000000000010;     //324pi/512
   m_cos[324]  =  15'b111111101011111;     //324pi/512
   m_sin[325]  =  15'b110000000000010;     //325pi/512
   m_cos[325]  =  15'b111111100110111;     //325pi/512
   m_sin[326]  =  15'b110000000000100;     //326pi/512
   m_cos[326]  =  15'b111111100001111;     //326pi/512
   m_sin[327]  =  15'b110000000000101;     //327pi/512
   m_cos[327]  =  15'b111111011100111;     //327pi/512
   m_sin[328]  =  15'b110000000000110;     //328pi/512
   m_cos[328]  =  15'b111111010111110;     //328pi/512
   m_sin[329]  =  15'b110000000001000;     //329pi/512
   m_cos[329]  =  15'b111111010010110;     //329pi/512
   m_sin[330]  =  15'b110000000001010;     //330pi/512
   m_cos[330]  =  15'b111111001101110;     //330pi/512
   m_sin[331]  =  15'b110000000001100;     //331pi/512
   m_cos[331]  =  15'b111111001000110;     //331pi/512
   m_sin[332]  =  15'b110000000001110;     //332pi/512
   m_cos[332]  =  15'b111111000011110;     //332pi/512
   m_sin[333]  =  15'b110000000010001;     //333pi/512
   m_cos[333]  =  15'b111110111110110;     //333pi/512
   m_sin[334]  =  15'b110000000010011;     //334pi/512
   m_cos[334]  =  15'b111110111001101;     //334pi/512
   m_sin[335]  =  15'b110000000010110;     //335pi/512
   m_cos[335]  =  15'b111110110100101;     //335pi/512
   m_sin[336]  =  15'b110000000011001;     //336pi/512
   m_cos[336]  =  15'b111110101111101;     //336pi/512
   m_sin[337]  =  15'b110000000011101;     //337pi/512
   m_cos[337]  =  15'b111110101010101;     //337pi/512
   m_sin[338]  =  15'b110000000100000;     //338pi/512
   m_cos[338]  =  15'b111110100101101;     //338pi/512
   m_sin[339]  =  15'b110000000100100;     //339pi/512
   m_cos[339]  =  15'b111110100000101;     //339pi/512
   m_sin[340]  =  15'b110000000100111;     //340pi/512
   m_cos[340]  =  15'b111110011011101;     //340pi/512
   m_sin[341]  =  15'b110000000101011;     //341pi/512
   m_cos[341]  =  15'b111110010110101;     //341pi/512
   m_sin[342]  =  15'b110000000110000;     //342pi/512
   m_cos[342]  =  15'b111110010001101;     //342pi/512
   m_sin[343]  =  15'b110000000110100;     //343pi/512
   m_cos[343]  =  15'b111110001100101;     //343pi/512
   m_sin[344]  =  15'b110000000111001;     //344pi/512
   m_cos[344]  =  15'b111110000111101;     //344pi/512
   m_sin[345]  =  15'b110000000111110;     //345pi/512
   m_cos[345]  =  15'b111110000010101;     //345pi/512
   m_sin[346]  =  15'b110000001000011;     //346pi/512
   m_cos[346]  =  15'b111101111101101;     //346pi/512
   m_sin[347]  =  15'b110000001001000;     //347pi/512
   m_cos[347]  =  15'b111101111000101;     //347pi/512
   m_sin[348]  =  15'b110000001001101;     //348pi/512
   m_cos[348]  =  15'b111101110011110;     //348pi/512
   m_sin[349]  =  15'b110000001010011;     //349pi/512
   m_cos[349]  =  15'b111101101110110;     //349pi/512
   m_sin[350]  =  15'b110000001011001;     //350pi/512
   m_cos[350]  =  15'b111101101001110;     //350pi/512
   m_sin[351]  =  15'b110000001011111;     //351pi/512
   m_cos[351]  =  15'b111101100100110;     //351pi/512
   m_sin[352]  =  15'b110000001100101;     //352pi/512
   m_cos[352]  =  15'b111101011111110;     //352pi/512
   m_sin[353]  =  15'b110000001101011;     //353pi/512
   m_cos[353]  =  15'b111101011010111;     //353pi/512
   m_sin[354]  =  15'b110000001110010;     //354pi/512
   m_cos[354]  =  15'b111101010101111;     //354pi/512
   m_sin[355]  =  15'b110000001111001;     //355pi/512
   m_cos[355]  =  15'b111101010000111;     //355pi/512
   m_sin[356]  =  15'b110000010000000;     //356pi/512
   m_cos[356]  =  15'b111101001100000;     //356pi/512
   m_sin[357]  =  15'b110000010000111;     //357pi/512
   m_cos[357]  =  15'b111101000111000;     //357pi/512
   m_sin[358]  =  15'b110000010001110;     //358pi/512
   m_cos[358]  =  15'b111101000010001;     //358pi/512
   m_sin[359]  =  15'b110000010010110;     //359pi/512
   m_cos[359]  =  15'b111100111101001;     //359pi/512
   m_sin[360]  =  15'b110000010011101;     //360pi/512
   m_cos[360]  =  15'b111100111000010;     //360pi/512
   m_sin[361]  =  15'b110000010100101;     //361pi/512
   m_cos[361]  =  15'b111100110011010;     //361pi/512
   m_sin[362]  =  15'b110000010101101;     //362pi/512
   m_cos[362]  =  15'b111100101110011;     //362pi/512
   m_sin[363]  =  15'b110000010110110;     //363pi/512
   m_cos[363]  =  15'b111100101001100;     //363pi/512
   m_sin[364]  =  15'b110000010111110;     //364pi/512
   m_cos[364]  =  15'b111100100100100;     //364pi/512
   m_sin[365]  =  15'b110000011000111;     //365pi/512
   m_cos[365]  =  15'b111100011111101;     //365pi/512
   m_sin[366]  =  15'b110000011010000;     //366pi/512
   m_cos[366]  =  15'b111100011010110;     //366pi/512
   m_sin[367]  =  15'b110000011011001;     //367pi/512
   m_cos[367]  =  15'b111100010101111;     //367pi/512
   m_sin[368]  =  15'b110000011100010;     //368pi/512
   m_cos[368]  =  15'b111100010001000;     //368pi/512
   m_sin[369]  =  15'b110000011101100;     //369pi/512
   m_cos[369]  =  15'b111100001100001;     //369pi/512
   m_sin[370]  =  15'b110000011110110;     //370pi/512
   m_cos[370]  =  15'b111100000111010;     //370pi/512
   m_sin[371]  =  15'b110000011111111;     //371pi/512
   m_cos[371]  =  15'b111100000010011;     //371pi/512
   m_sin[372]  =  15'b110000100001001;     //372pi/512
   m_cos[372]  =  15'b111011111101100;     //372pi/512
   m_sin[373]  =  15'b110000100010100;     //373pi/512
   m_cos[373]  =  15'b111011111000101;     //373pi/512
   m_sin[374]  =  15'b110000100011110;     //374pi/512
   m_cos[374]  =  15'b111011110011110;     //374pi/512
   m_sin[375]  =  15'b110000100101001;     //375pi/512
   m_cos[375]  =  15'b111011101110111;     //375pi/512
   m_sin[376]  =  15'b110000100110100;     //376pi/512
   m_cos[376]  =  15'b111011101010000;     //376pi/512
   m_sin[377]  =  15'b110000100111111;     //377pi/512
   m_cos[377]  =  15'b111011100101010;     //377pi/512
   m_sin[378]  =  15'b110000101001010;     //378pi/512
   m_cos[378]  =  15'b111011100000011;     //378pi/512
   m_sin[379]  =  15'b110000101010101;     //379pi/512
   m_cos[379]  =  15'b111011011011100;     //379pi/512
   m_sin[380]  =  15'b110000101100001;     //380pi/512
   m_cos[380]  =  15'b111011010110110;     //380pi/512
   m_sin[381]  =  15'b110000101101101;     //381pi/512
   m_cos[381]  =  15'b111011010010000;     //381pi/512
   m_sin[382]  =  15'b110000101111000;     //382pi/512
   m_cos[382]  =  15'b111011001101001;     //382pi/512
   m_sin[383]  =  15'b110000110000101;     //383pi/512
   m_cos[383]  =  15'b111011001000011;     //383pi/512
   m_sin[384]  =  15'b110000110010001;     //384pi/512
   m_cos[384]  =  15'b111011000011101;     //384pi/512
   m_sin[385]  =  15'b110000110011101;     //385pi/512
   m_cos[385]  =  15'b111010111110110;     //385pi/512
   m_sin[386]  =  15'b110000110101010;     //386pi/512
   m_cos[386]  =  15'b111010111010000;     //386pi/512
   m_sin[387]  =  15'b110000110110111;     //387pi/512
   m_cos[387]  =  15'b111010110101010;     //387pi/512
   m_sin[388]  =  15'b110000111000100;     //388pi/512
   m_cos[388]  =  15'b111010110000100;     //388pi/512
   m_sin[389]  =  15'b110000111010001;     //389pi/512
   m_cos[389]  =  15'b111010101011110;     //389pi/512
   m_sin[390]  =  15'b110000111011111;     //390pi/512
   m_cos[390]  =  15'b111010100111000;     //390pi/512
   m_sin[391]  =  15'b110000111101101;     //391pi/512
   m_cos[391]  =  15'b111010100010010;     //391pi/512
   m_sin[392]  =  15'b110000111111010;     //392pi/512
   m_cos[392]  =  15'b111010011101101;     //392pi/512
   m_sin[393]  =  15'b110001000001000;     //393pi/512
   m_cos[393]  =  15'b111010011000111;     //393pi/512
   m_sin[394]  =  15'b110001000010111;     //394pi/512
   m_cos[394]  =  15'b111010010100001;     //394pi/512
   m_sin[395]  =  15'b110001000100101;     //395pi/512
   m_cos[395]  =  15'b111010001111100;     //395pi/512
   m_sin[396]  =  15'b110001000110011;     //396pi/512
   m_cos[396]  =  15'b111010001010110;     //396pi/512
   m_sin[397]  =  15'b110001001000010;     //397pi/512
   m_cos[397]  =  15'b111010000110001;     //397pi/512
   m_sin[398]  =  15'b110001001010001;     //398pi/512
   m_cos[398]  =  15'b111010000001100;     //398pi/512
   m_sin[399]  =  15'b110001001100000;     //399pi/512
   m_cos[399]  =  15'b111001111100110;     //399pi/512
   m_sin[400]  =  15'b110001001110000;     //400pi/512
   m_cos[400]  =  15'b111001111000001;     //400pi/512
   m_sin[401]  =  15'b110001001111111;     //401pi/512
   m_cos[401]  =  15'b111001110011100;     //401pi/512
   m_sin[402]  =  15'b110001010001111;     //402pi/512
   m_cos[402]  =  15'b111001101110111;     //402pi/512
   m_sin[403]  =  15'b110001010011111;     //403pi/512
   m_cos[403]  =  15'b111001101010010;     //403pi/512
   m_sin[404]  =  15'b110001010101111;     //404pi/512
   m_cos[404]  =  15'b111001100101101;     //404pi/512
   m_sin[405]  =  15'b110001010111111;     //405pi/512
   m_cos[405]  =  15'b111001100001000;     //405pi/512
   m_sin[406]  =  15'b110001011001111;     //406pi/512
   m_cos[406]  =  15'b111001011100100;     //406pi/512
   m_sin[407]  =  15'b110001011100000;     //407pi/512
   m_cos[407]  =  15'b111001010111111;     //407pi/512
   m_sin[408]  =  15'b110001011110000;     //408pi/512
   m_cos[408]  =  15'b111001010011010;     //408pi/512
   m_sin[409]  =  15'b110001100000001;     //409pi/512
   m_cos[409]  =  15'b111001001110110;     //409pi/512
   m_sin[410]  =  15'b110001100010011;     //410pi/512
   m_cos[410]  =  15'b111001001010001;     //410pi/512
   m_sin[411]  =  15'b110001100100100;     //411pi/512
   m_cos[411]  =  15'b111001000101101;     //411pi/512
   m_sin[412]  =  15'b110001100110101;     //412pi/512
   m_cos[412]  =  15'b111001000001001;     //412pi/512
   m_sin[413]  =  15'b110001101000111;     //413pi/512
   m_cos[413]  =  15'b111000111100101;     //413pi/512
   m_sin[414]  =  15'b110001101011001;     //414pi/512
   m_cos[414]  =  15'b111000111000001;     //414pi/512
   m_sin[415]  =  15'b110001101101011;     //415pi/512
   m_cos[415]  =  15'b111000110011101;     //415pi/512
   m_sin[416]  =  15'b110001101111101;     //416pi/512
   m_cos[416]  =  15'b111000101111001;     //416pi/512
   m_sin[417]  =  15'b110001110001111;     //417pi/512
   m_cos[417]  =  15'b111000101010101;     //417pi/512
   m_sin[418]  =  15'b110001110100010;     //418pi/512
   m_cos[418]  =  15'b111000100110001;     //418pi/512
   m_sin[419]  =  15'b110001110110100;     //419pi/512
   m_cos[419]  =  15'b111000100001110;     //419pi/512
   m_sin[420]  =  15'b110001111000111;     //420pi/512
   m_cos[420]  =  15'b111000011101010;     //420pi/512
   m_sin[421]  =  15'b110001111011010;     //421pi/512
   m_cos[421]  =  15'b111000011000111;     //421pi/512
   m_sin[422]  =  15'b110001111101110;     //422pi/512
   m_cos[422]  =  15'b111000010100100;     //422pi/512
   m_sin[423]  =  15'b110010000000001;     //423pi/512
   m_cos[423]  =  15'b111000010000000;     //423pi/512
   m_sin[424]  =  15'b110010000010101;     //424pi/512
   m_cos[424]  =  15'b111000001011101;     //424pi/512
   m_sin[425]  =  15'b110010000101000;     //425pi/512
   m_cos[425]  =  15'b111000000111010;     //425pi/512
   m_sin[426]  =  15'b110010000111100;     //426pi/512
   m_cos[426]  =  15'b111000000010111;     //426pi/512
   m_sin[427]  =  15'b110010001010000;     //427pi/512
   m_cos[427]  =  15'b110111111110100;     //427pi/512
   m_sin[428]  =  15'b110010001100100;     //428pi/512
   m_cos[428]  =  15'b110111111010010;     //428pi/512
   m_sin[429]  =  15'b110010001111001;     //429pi/512
   m_cos[429]  =  15'b110111110101111;     //429pi/512
   m_sin[430]  =  15'b110010010001101;     //430pi/512
   m_cos[430]  =  15'b110111110001100;     //430pi/512
   m_sin[431]  =  15'b110010010100010;     //431pi/512
   m_cos[431]  =  15'b110111101101010;     //431pi/512
   m_sin[432]  =  15'b110010010110111;     //432pi/512
   m_cos[432]  =  15'b110111101001000;     //432pi/512
   m_sin[433]  =  15'b110010011001100;     //433pi/512
   m_cos[433]  =  15'b110111100100101;     //433pi/512
   m_sin[434]  =  15'b110010011100010;     //434pi/512
   m_cos[434]  =  15'b110111100000011;     //434pi/512
   m_sin[435]  =  15'b110010011110111;     //435pi/512
   m_cos[435]  =  15'b110111011100001;     //435pi/512
   m_sin[436]  =  15'b110010100001101;     //436pi/512
   m_cos[436]  =  15'b110111010111111;     //436pi/512
   m_sin[437]  =  15'b110010100100010;     //437pi/512
   m_cos[437]  =  15'b110111010011110;     //437pi/512
   m_sin[438]  =  15'b110010100111000;     //438pi/512
   m_cos[438]  =  15'b110111001111100;     //438pi/512
   m_sin[439]  =  15'b110010101001110;     //439pi/512
   m_cos[439]  =  15'b110111001011010;     //439pi/512
   m_sin[440]  =  15'b110010101100101;     //440pi/512
   m_cos[440]  =  15'b110111000111001;     //440pi/512
   m_sin[441]  =  15'b110010101111011;     //441pi/512
   m_cos[441]  =  15'b110111000010111;     //441pi/512
   m_sin[442]  =  15'b110010110010010;     //442pi/512
   m_cos[442]  =  15'b110110111110110;     //442pi/512
   m_sin[443]  =  15'b110010110101000;     //443pi/512
   m_cos[443]  =  15'b110110111010101;     //443pi/512
   m_sin[444]  =  15'b110010110111111;     //444pi/512
   m_cos[444]  =  15'b110110110110100;     //444pi/512
   m_sin[445]  =  15'b110010111010110;     //445pi/512
   m_cos[445]  =  15'b110110110010011;     //445pi/512
   m_sin[446]  =  15'b110010111101110;     //446pi/512
   m_cos[446]  =  15'b110110101110010;     //446pi/512
   m_sin[447]  =  15'b110011000000101;     //447pi/512
   m_cos[447]  =  15'b110110101010001;     //447pi/512
   m_sin[448]  =  15'b110011000011101;     //448pi/512
   m_cos[448]  =  15'b110110100110001;     //448pi/512
   m_sin[449]  =  15'b110011000110100;     //449pi/512
   m_cos[449]  =  15'b110110100010000;     //449pi/512
   m_sin[450]  =  15'b110011001001100;     //450pi/512
   m_cos[450]  =  15'b110110011110000;     //450pi/512
   m_sin[451]  =  15'b110011001100100;     //451pi/512
   m_cos[451]  =  15'b110110011010000;     //451pi/512
   m_sin[452]  =  15'b110011001111100;     //452pi/512
   m_cos[452]  =  15'b110110010110000;     //452pi/512
   m_sin[453]  =  15'b110011010010101;     //453pi/512
   m_cos[453]  =  15'b110110010010000;     //453pi/512
   m_sin[454]  =  15'b110011010101101;     //454pi/512
   m_cos[454]  =  15'b110110001110000;     //454pi/512
   m_sin[455]  =  15'b110011011000110;     //455pi/512
   m_cos[455]  =  15'b110110001010000;     //455pi/512
   m_sin[456]  =  15'b110011011011111;     //456pi/512
   m_cos[456]  =  15'b110110000110000;     //456pi/512
   m_sin[457]  =  15'b110011011111000;     //457pi/512
   m_cos[457]  =  15'b110110000010001;     //457pi/512
   m_sin[458]  =  15'b110011100010001;     //458pi/512
   m_cos[458]  =  15'b110101111110001;     //458pi/512
   m_sin[459]  =  15'b110011100101010;     //459pi/512
   m_cos[459]  =  15'b110101111010010;     //459pi/512
   m_sin[460]  =  15'b110011101000011;     //460pi/512
   m_cos[460]  =  15'b110101110110011;     //460pi/512
   m_sin[461]  =  15'b110011101011101;     //461pi/512
   m_cos[461]  =  15'b110101110010100;     //461pi/512
   m_sin[462]  =  15'b110011101110111;     //462pi/512
   m_cos[462]  =  15'b110101101110101;     //462pi/512
   m_sin[463]  =  15'b110011110010001;     //463pi/512
   m_cos[463]  =  15'b110101101010110;     //463pi/512
   m_sin[464]  =  15'b110011110101011;     //464pi/512
   m_cos[464]  =  15'b110101100111000;     //464pi/512
   m_sin[465]  =  15'b110011111000101;     //465pi/512
   m_cos[465]  =  15'b110101100011001;     //465pi/512
   m_sin[466]  =  15'b110011111011111;     //466pi/512
   m_cos[466]  =  15'b110101011111011;     //466pi/512
   m_sin[467]  =  15'b110011111111010;     //467pi/512
   m_cos[467]  =  15'b110101011011101;     //467pi/512
   m_sin[468]  =  15'b110100000010100;     //468pi/512
   m_cos[468]  =  15'b110101010111110;     //468pi/512
   m_sin[469]  =  15'b110100000101111;     //469pi/512
   m_cos[469]  =  15'b110101010100000;     //469pi/512
   m_sin[470]  =  15'b110100001001010;     //470pi/512
   m_cos[470]  =  15'b110101010000011;     //470pi/512
   m_sin[471]  =  15'b110100001100101;     //471pi/512
   m_cos[471]  =  15'b110101001100101;     //471pi/512
   m_sin[472]  =  15'b110100010000000;     //472pi/512
   m_cos[472]  =  15'b110101001000111;     //472pi/512
   m_sin[473]  =  15'b110100010011100;     //473pi/512
   m_cos[473]  =  15'b110101000101010;     //473pi/512
   m_sin[474]  =  15'b110100010110111;     //474pi/512
   m_cos[474]  =  15'b110101000001100;     //474pi/512
   m_sin[475]  =  15'b110100011010011;     //475pi/512
   m_cos[475]  =  15'b110100111101111;     //475pi/512
   m_sin[476]  =  15'b110100011101111;     //476pi/512
   m_cos[476]  =  15'b110100111010010;     //476pi/512
   m_sin[477]  =  15'b110100100001011;     //477pi/512
   m_cos[477]  =  15'b110100110110101;     //477pi/512
   m_sin[478]  =  15'b110100100100111;     //478pi/512
   m_cos[478]  =  15'b110100110011001;     //478pi/512
   m_sin[479]  =  15'b110100101000011;     //479pi/512
   m_cos[479]  =  15'b110100101111100;     //479pi/512
   m_sin[480]  =  15'b110100101011111;     //480pi/512
   m_cos[480]  =  15'b110100101011111;     //480pi/512
   m_sin[481]  =  15'b110100101111100;     //481pi/512
   m_cos[481]  =  15'b110100101000011;     //481pi/512
   m_sin[482]  =  15'b110100110011001;     //482pi/512
   m_cos[482]  =  15'b110100100100111;     //482pi/512
   m_sin[483]  =  15'b110100110110101;     //483pi/512
   m_cos[483]  =  15'b110100100001011;     //483pi/512
   m_sin[484]  =  15'b110100111010010;     //484pi/512
   m_cos[484]  =  15'b110100011101111;     //484pi/512
   m_sin[485]  =  15'b110100111101111;     //485pi/512
   m_cos[485]  =  15'b110100011010011;     //485pi/512
   m_sin[486]  =  15'b110101000001100;     //486pi/512
   m_cos[486]  =  15'b110100010110111;     //486pi/512
   m_sin[487]  =  15'b110101000101010;     //487pi/512
   m_cos[487]  =  15'b110100010011100;     //487pi/512
   m_sin[488]  =  15'b110101001000111;     //488pi/512
   m_cos[488]  =  15'b110100010000000;     //488pi/512
   m_sin[489]  =  15'b110101001100101;     //489pi/512
   m_cos[489]  =  15'b110100001100101;     //489pi/512
   m_sin[490]  =  15'b110101010000011;     //490pi/512
   m_cos[490]  =  15'b110100001001010;     //490pi/512
   m_sin[491]  =  15'b110101010100000;     //491pi/512
   m_cos[491]  =  15'b110100000101111;     //491pi/512
   m_sin[492]  =  15'b110101010111110;     //492pi/512
   m_cos[492]  =  15'b110100000010100;     //492pi/512
   m_sin[493]  =  15'b110101011011101;     //493pi/512
   m_cos[493]  =  15'b110011111111010;     //493pi/512
   m_sin[494]  =  15'b110101011111011;     //494pi/512
   m_cos[494]  =  15'b110011111011111;     //494pi/512
   m_sin[495]  =  15'b110101100011001;     //495pi/512
   m_cos[495]  =  15'b110011111000101;     //495pi/512
   m_sin[496]  =  15'b110101100111000;     //496pi/512
   m_cos[496]  =  15'b110011110101011;     //496pi/512
   m_sin[497]  =  15'b110101101010110;     //497pi/512
   m_cos[497]  =  15'b110011110010001;     //497pi/512
   m_sin[498]  =  15'b110101101110101;     //498pi/512
   m_cos[498]  =  15'b110011101110111;     //498pi/512
   m_sin[499]  =  15'b110101110010100;     //499pi/512
   m_cos[499]  =  15'b110011101011101;     //499pi/512
   m_sin[500]  =  15'b110101110110011;     //500pi/512
   m_cos[500]  =  15'b110011101000011;     //500pi/512
   m_sin[501]  =  15'b110101111010010;     //501pi/512
   m_cos[501]  =  15'b110011100101010;     //501pi/512
   m_sin[502]  =  15'b110101111110001;     //502pi/512
   m_cos[502]  =  15'b110011100010001;     //502pi/512
   m_sin[503]  =  15'b110110000010001;     //503pi/512
   m_cos[503]  =  15'b110011011111000;     //503pi/512
   m_sin[504]  =  15'b110110000110000;     //504pi/512
   m_cos[504]  =  15'b110011011011111;     //504pi/512
   m_sin[505]  =  15'b110110001010000;     //505pi/512
   m_cos[505]  =  15'b110011011000110;     //505pi/512
   m_sin[506]  =  15'b110110001110000;     //506pi/512
   m_cos[506]  =  15'b110011010101101;     //506pi/512
   m_sin[507]  =  15'b110110010010000;     //507pi/512
   m_cos[507]  =  15'b110011010010101;     //507pi/512
   m_sin[508]  =  15'b110110010110000;     //508pi/512
   m_cos[508]  =  15'b110011001111100;     //508pi/512
   m_sin[509]  =  15'b110110011010000;     //509pi/512
   m_cos[509]  =  15'b110011001100100;     //509pi/512
   m_sin[510]  =  15'b110110011110000;     //510pi/512
   m_cos[510]  =  15'b110011001001100;     //510pi/512
   m_sin[511]  =  15'b110110100010000;     //511pi/512
   m_cos[511]  =  15'b110011000110100;     //511pi/512
end
endmodule
