module  M_TWIDLE_10_bit #(parameter SIZE =10, word_length_tw = 10) (
    input            clk,
    input            en_rd, 
    input   [10:0]   rd_ptr_angle,
    input            en_modf, 

    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );


reg signed [word_length_tw-1:0]  cos  [511:0];
reg signed [word_length_tw-1:0]  sin  [511:0];

reg signed [word_length_tw-1:0]  m_cos  [511:0];
reg signed [word_length_tw-1:0]  m_sin  [511:0];

reg signed [word_length_tw-1:0]  cos_temp;
reg signed [word_length_tw-1:0]  sin_temp;

reg signed [word_length_tw-1:0]  m_cos_temp;
reg signed [word_length_tw-1:0]  m_sin_temp;


//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & ~ en_modf ) begin
                  cos_temp           <= cos   [rd_ptr_angle];
                  sin_temp           <= sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & en_modf ) begin
                  m_cos_temp           <= m_cos   [rd_ptr_angle];
                  m_sin_temp           <= m_sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(*) begin 
             if (en_modf ) begin
                  cos_data           <= m_cos_temp;
                  sin_data           <= m_sin_temp;
             end else begin
                  cos_data           <= cos_temp;
                  sin_data           <= sin_temp;
             end
        end
//----------------------------------------------------------------------------------------
initial begin
   sin[0]  =  10'b0000000000;     //0pi/512
   cos[0]  =  10'b0100000000;     //0pi/512
   sin[1]  =  10'b1111111110;     //1pi/512
   cos[1]  =  10'b0011111111;     //1pi/512
   sin[2]  =  10'b1111111101;     //2pi/512
   cos[2]  =  10'b0011111111;     //2pi/512
   sin[3]  =  10'b1111111011;     //3pi/512
   cos[3]  =  10'b0011111111;     //3pi/512
   sin[4]  =  10'b1111111010;     //4pi/512
   cos[4]  =  10'b0011111111;     //4pi/512
   sin[5]  =  10'b1111111000;     //5pi/512
   cos[5]  =  10'b0011111111;     //5pi/512
   sin[6]  =  10'b1111110111;     //6pi/512
   cos[6]  =  10'b0011111111;     //6pi/512
   sin[7]  =  10'b1111110101;     //7pi/512
   cos[7]  =  10'b0011111111;     //7pi/512
   sin[8]  =  10'b1111110011;     //8pi/512
   cos[8]  =  10'b0011111111;     //8pi/512
   sin[9]  =  10'b1111110010;     //9pi/512
   cos[9]  =  10'b0011111111;     //9pi/512
   sin[10]  =  10'b1111110000;     //10pi/512
   cos[10]  =  10'b0011111111;     //10pi/512
   sin[11]  =  10'b1111101111;     //11pi/512
   cos[11]  =  10'b0011111111;     //11pi/512
   sin[12]  =  10'b1111101101;     //12pi/512
   cos[12]  =  10'b0011111111;     //12pi/512
   sin[13]  =  10'b1111101100;     //13pi/512
   cos[13]  =  10'b0011111111;     //13pi/512
   sin[14]  =  10'b1111101010;     //14pi/512
   cos[14]  =  10'b0011111111;     //14pi/512
   sin[15]  =  10'b1111101000;     //15pi/512
   cos[15]  =  10'b0011111110;     //15pi/512
   sin[16]  =  10'b1111100111;     //16pi/512
   cos[16]  =  10'b0011111110;     //16pi/512
   sin[17]  =  10'b1111100101;     //17pi/512
   cos[17]  =  10'b0011111110;     //17pi/512
   sin[18]  =  10'b1111100100;     //18pi/512
   cos[18]  =  10'b0011111110;     //18pi/512
   sin[19]  =  10'b1111100010;     //19pi/512
   cos[19]  =  10'b0011111110;     //19pi/512
   sin[20]  =  10'b1111100001;     //20pi/512
   cos[20]  =  10'b0011111110;     //20pi/512
   sin[21]  =  10'b1111011111;     //21pi/512
   cos[21]  =  10'b0011111101;     //21pi/512
   sin[22]  =  10'b1111011110;     //22pi/512
   cos[22]  =  10'b0011111101;     //22pi/512
   sin[23]  =  10'b1111011100;     //23pi/512
   cos[23]  =  10'b0011111101;     //23pi/512
   sin[24]  =  10'b1111011010;     //24pi/512
   cos[24]  =  10'b0011111101;     //24pi/512
   sin[25]  =  10'b1111011001;     //25pi/512
   cos[25]  =  10'b0011111100;     //25pi/512
   sin[26]  =  10'b1111010111;     //26pi/512
   cos[26]  =  10'b0011111100;     //26pi/512
   sin[27]  =  10'b1111010110;     //27pi/512
   cos[27]  =  10'b0011111100;     //27pi/512
   sin[28]  =  10'b1111010100;     //28pi/512
   cos[28]  =  10'b0011111100;     //28pi/512
   sin[29]  =  10'b1111010011;     //29pi/512
   cos[29]  =  10'b0011111011;     //29pi/512
   sin[30]  =  10'b1111010001;     //30pi/512
   cos[30]  =  10'b0011111011;     //30pi/512
   sin[31]  =  10'b1111010000;     //31pi/512
   cos[31]  =  10'b0011111011;     //31pi/512
   sin[32]  =  10'b1111001110;     //32pi/512
   cos[32]  =  10'b0011111011;     //32pi/512
   sin[33]  =  10'b1111001101;     //33pi/512
   cos[33]  =  10'b0011111010;     //33pi/512
   sin[34]  =  10'b1111001011;     //34pi/512
   cos[34]  =  10'b0011111010;     //34pi/512
   sin[35]  =  10'b1111001001;     //35pi/512
   cos[35]  =  10'b0011111010;     //35pi/512
   sin[36]  =  10'b1111001000;     //36pi/512
   cos[36]  =  10'b0011111001;     //36pi/512
   sin[37]  =  10'b1111000110;     //37pi/512
   cos[37]  =  10'b0011111001;     //37pi/512
   sin[38]  =  10'b1111000101;     //38pi/512
   cos[38]  =  10'b0011111001;     //38pi/512
   sin[39]  =  10'b1111000011;     //39pi/512
   cos[39]  =  10'b0011111000;     //39pi/512
   sin[40]  =  10'b1111000010;     //40pi/512
   cos[40]  =  10'b0011111000;     //40pi/512
   sin[41]  =  10'b1111000000;     //41pi/512
   cos[41]  =  10'b0011110111;     //41pi/512
   sin[42]  =  10'b1110111111;     //42pi/512
   cos[42]  =  10'b0011110111;     //42pi/512
   sin[43]  =  10'b1110111101;     //43pi/512
   cos[43]  =  10'b0011110111;     //43pi/512
   sin[44]  =  10'b1110111100;     //44pi/512
   cos[44]  =  10'b0011110110;     //44pi/512
   sin[45]  =  10'b1110111010;     //45pi/512
   cos[45]  =  10'b0011110110;     //45pi/512
   sin[46]  =  10'b1110111001;     //46pi/512
   cos[46]  =  10'b0011110101;     //46pi/512
   sin[47]  =  10'b1110110111;     //47pi/512
   cos[47]  =  10'b0011110101;     //47pi/512
   sin[48]  =  10'b1110110110;     //48pi/512
   cos[48]  =  10'b0011110100;     //48pi/512
   sin[49]  =  10'b1110110100;     //49pi/512
   cos[49]  =  10'b0011110100;     //49pi/512
   sin[50]  =  10'b1110110011;     //50pi/512
   cos[50]  =  10'b0011110100;     //50pi/512
   sin[51]  =  10'b1110110001;     //51pi/512
   cos[51]  =  10'b0011110011;     //51pi/512
   sin[52]  =  10'b1110110000;     //52pi/512
   cos[52]  =  10'b0011110011;     //52pi/512
   sin[53]  =  10'b1110101110;     //53pi/512
   cos[53]  =  10'b0011110010;     //53pi/512
   sin[54]  =  10'b1110101101;     //54pi/512
   cos[54]  =  10'b0011110010;     //54pi/512
   sin[55]  =  10'b1110101011;     //55pi/512
   cos[55]  =  10'b0011110001;     //55pi/512
   sin[56]  =  10'b1110101010;     //56pi/512
   cos[56]  =  10'b0011110001;     //56pi/512
   sin[57]  =  10'b1110101000;     //57pi/512
   cos[57]  =  10'b0011110000;     //57pi/512
   sin[58]  =  10'b1110100111;     //58pi/512
   cos[58]  =  10'b0011101111;     //58pi/512
   sin[59]  =  10'b1110100101;     //59pi/512
   cos[59]  =  10'b0011101111;     //59pi/512
   sin[60]  =  10'b1110100100;     //60pi/512
   cos[60]  =  10'b0011101110;     //60pi/512
   sin[61]  =  10'b1110100010;     //61pi/512
   cos[61]  =  10'b0011101110;     //61pi/512
   sin[62]  =  10'b1110100001;     //62pi/512
   cos[62]  =  10'b0011101101;     //62pi/512
   sin[63]  =  10'b1110011111;     //63pi/512
   cos[63]  =  10'b0011101101;     //63pi/512
   sin[64]  =  10'b1110011110;     //64pi/512
   cos[64]  =  10'b0011101100;     //64pi/512
   sin[65]  =  10'b1110011101;     //65pi/512
   cos[65]  =  10'b0011101011;     //65pi/512
   sin[66]  =  10'b1110011011;     //66pi/512
   cos[66]  =  10'b0011101011;     //66pi/512
   sin[67]  =  10'b1110011010;     //67pi/512
   cos[67]  =  10'b0011101010;     //67pi/512
   sin[68]  =  10'b1110011000;     //68pi/512
   cos[68]  =  10'b0011101010;     //68pi/512
   sin[69]  =  10'b1110010111;     //69pi/512
   cos[69]  =  10'b0011101001;     //69pi/512
   sin[70]  =  10'b1110010101;     //70pi/512
   cos[70]  =  10'b0011101000;     //70pi/512
   sin[71]  =  10'b1110010100;     //71pi/512
   cos[71]  =  10'b0011101000;     //71pi/512
   sin[72]  =  10'b1110010011;     //72pi/512
   cos[72]  =  10'b0011100111;     //72pi/512
   sin[73]  =  10'b1110010001;     //73pi/512
   cos[73]  =  10'b0011100110;     //73pi/512
   sin[74]  =  10'b1110010000;     //74pi/512
   cos[74]  =  10'b0011100110;     //74pi/512
   sin[75]  =  10'b1110001110;     //75pi/512
   cos[75]  =  10'b0011100101;     //75pi/512
   sin[76]  =  10'b1110001101;     //76pi/512
   cos[76]  =  10'b0011100100;     //76pi/512
   sin[77]  =  10'b1110001011;     //77pi/512
   cos[77]  =  10'b0011100011;     //77pi/512
   sin[78]  =  10'b1110001010;     //78pi/512
   cos[78]  =  10'b0011100011;     //78pi/512
   sin[79]  =  10'b1110001001;     //79pi/512
   cos[79]  =  10'b0011100010;     //79pi/512
   sin[80]  =  10'b1110000111;     //80pi/512
   cos[80]  =  10'b0011100001;     //80pi/512
   sin[81]  =  10'b1110000110;     //81pi/512
   cos[81]  =  10'b0011100001;     //81pi/512
   sin[82]  =  10'b1110000101;     //82pi/512
   cos[82]  =  10'b0011100000;     //82pi/512
   sin[83]  =  10'b1110000011;     //83pi/512
   cos[83]  =  10'b0011011111;     //83pi/512
   sin[84]  =  10'b1110000010;     //84pi/512
   cos[84]  =  10'b0011011110;     //84pi/512
   sin[85]  =  10'b1110000000;     //85pi/512
   cos[85]  =  10'b0011011101;     //85pi/512
   sin[86]  =  10'b1101111111;     //86pi/512
   cos[86]  =  10'b0011011101;     //86pi/512
   sin[87]  =  10'b1101111110;     //87pi/512
   cos[87]  =  10'b0011011100;     //87pi/512
   sin[88]  =  10'b1101111100;     //88pi/512
   cos[88]  =  10'b0011011011;     //88pi/512
   sin[89]  =  10'b1101111011;     //89pi/512
   cos[89]  =  10'b0011011010;     //89pi/512
   sin[90]  =  10'b1101111010;     //90pi/512
   cos[90]  =  10'b0011011001;     //90pi/512
   sin[91]  =  10'b1101111000;     //91pi/512
   cos[91]  =  10'b0011011001;     //91pi/512
   sin[92]  =  10'b1101110111;     //92pi/512
   cos[92]  =  10'b0011011000;     //92pi/512
   sin[93]  =  10'b1101110110;     //93pi/512
   cos[93]  =  10'b0011010111;     //93pi/512
   sin[94]  =  10'b1101110100;     //94pi/512
   cos[94]  =  10'b0011010110;     //94pi/512
   sin[95]  =  10'b1101110011;     //95pi/512
   cos[95]  =  10'b0011010101;     //95pi/512
   sin[96]  =  10'b1101110010;     //96pi/512
   cos[96]  =  10'b0011010100;     //96pi/512
   sin[97]  =  10'b1101110000;     //97pi/512
   cos[97]  =  10'b0011010011;     //97pi/512
   sin[98]  =  10'b1101101111;     //98pi/512
   cos[98]  =  10'b0011010011;     //98pi/512
   sin[99]  =  10'b1101101110;     //99pi/512
   cos[99]  =  10'b0011010010;     //99pi/512
   sin[100]  =  10'b1101101101;     //100pi/512
   cos[100]  =  10'b0011010001;     //100pi/512
   sin[101]  =  10'b1101101011;     //101pi/512
   cos[101]  =  10'b0011010000;     //101pi/512
   sin[102]  =  10'b1101101010;     //102pi/512
   cos[102]  =  10'b0011001111;     //102pi/512
   sin[103]  =  10'b1101101001;     //103pi/512
   cos[103]  =  10'b0011001110;     //103pi/512
   sin[104]  =  10'b1101101000;     //104pi/512
   cos[104]  =  10'b0011001101;     //104pi/512
   sin[105]  =  10'b1101100110;     //105pi/512
   cos[105]  =  10'b0011001100;     //105pi/512
   sin[106]  =  10'b1101100101;     //106pi/512
   cos[106]  =  10'b0011001011;     //106pi/512
   sin[107]  =  10'b1101100100;     //107pi/512
   cos[107]  =  10'b0011001010;     //107pi/512
   sin[108]  =  10'b1101100011;     //108pi/512
   cos[108]  =  10'b0011001001;     //108pi/512
   sin[109]  =  10'b1101100001;     //109pi/512
   cos[109]  =  10'b0011001000;     //109pi/512
   sin[110]  =  10'b1101100000;     //110pi/512
   cos[110]  =  10'b0011000111;     //110pi/512
   sin[111]  =  10'b1101011111;     //111pi/512
   cos[111]  =  10'b0011000110;     //111pi/512
   sin[112]  =  10'b1101011110;     //112pi/512
   cos[112]  =  10'b0011000101;     //112pi/512
   sin[113]  =  10'b1101011100;     //113pi/512
   cos[113]  =  10'b0011000100;     //113pi/512
   sin[114]  =  10'b1101011011;     //114pi/512
   cos[114]  =  10'b0011000011;     //114pi/512
   sin[115]  =  10'b1101011010;     //115pi/512
   cos[115]  =  10'b0011000010;     //115pi/512
   sin[116]  =  10'b1101011001;     //116pi/512
   cos[116]  =  10'b0011000001;     //116pi/512
   sin[117]  =  10'b1101011000;     //117pi/512
   cos[117]  =  10'b0011000000;     //117pi/512
   sin[118]  =  10'b1101010110;     //118pi/512
   cos[118]  =  10'b0010111111;     //118pi/512
   sin[119]  =  10'b1101010101;     //119pi/512
   cos[119]  =  10'b0010111110;     //119pi/512
   sin[120]  =  10'b1101010100;     //120pi/512
   cos[120]  =  10'b0010111101;     //120pi/512
   sin[121]  =  10'b1101010011;     //121pi/512
   cos[121]  =  10'b0010111100;     //121pi/512
   sin[122]  =  10'b1101010010;     //122pi/512
   cos[122]  =  10'b0010111011;     //122pi/512
   sin[123]  =  10'b1101010001;     //123pi/512
   cos[123]  =  10'b0010111010;     //123pi/512
   sin[124]  =  10'b1101001111;     //124pi/512
   cos[124]  =  10'b0010111001;     //124pi/512
   sin[125]  =  10'b1101001110;     //125pi/512
   cos[125]  =  10'b0010111000;     //125pi/512
   sin[126]  =  10'b1101001101;     //126pi/512
   cos[126]  =  10'b0010110111;     //126pi/512
   sin[127]  =  10'b1101001100;     //127pi/512
   cos[127]  =  10'b0010110110;     //127pi/512
   sin[128]  =  10'b1101001011;     //128pi/512
   cos[128]  =  10'b0010110101;     //128pi/512
   sin[129]  =  10'b1101001010;     //129pi/512
   cos[129]  =  10'b0010110011;     //129pi/512
   sin[130]  =  10'b1101001001;     //130pi/512
   cos[130]  =  10'b0010110010;     //130pi/512
   sin[131]  =  10'b1101001000;     //131pi/512
   cos[131]  =  10'b0010110001;     //131pi/512
   sin[132]  =  10'b1101000111;     //132pi/512
   cos[132]  =  10'b0010110000;     //132pi/512
   sin[133]  =  10'b1101000110;     //133pi/512
   cos[133]  =  10'b0010101111;     //133pi/512
   sin[134]  =  10'b1101000100;     //134pi/512
   cos[134]  =  10'b0010101110;     //134pi/512
   sin[135]  =  10'b1101000011;     //135pi/512
   cos[135]  =  10'b0010101101;     //135pi/512
   sin[136]  =  10'b1101000010;     //136pi/512
   cos[136]  =  10'b0010101011;     //136pi/512
   sin[137]  =  10'b1101000001;     //137pi/512
   cos[137]  =  10'b0010101010;     //137pi/512
   sin[138]  =  10'b1101000000;     //138pi/512
   cos[138]  =  10'b0010101001;     //138pi/512
   sin[139]  =  10'b1100111111;     //139pi/512
   cos[139]  =  10'b0010101000;     //139pi/512
   sin[140]  =  10'b1100111110;     //140pi/512
   cos[140]  =  10'b0010100111;     //140pi/512
   sin[141]  =  10'b1100111101;     //141pi/512
   cos[141]  =  10'b0010100110;     //141pi/512
   sin[142]  =  10'b1100111100;     //142pi/512
   cos[142]  =  10'b0010100100;     //142pi/512
   sin[143]  =  10'b1100111011;     //143pi/512
   cos[143]  =  10'b0010100011;     //143pi/512
   sin[144]  =  10'b1100111010;     //144pi/512
   cos[144]  =  10'b0010100010;     //144pi/512
   sin[145]  =  10'b1100111001;     //145pi/512
   cos[145]  =  10'b0010100001;     //145pi/512
   sin[146]  =  10'b1100111000;     //146pi/512
   cos[146]  =  10'b0010011111;     //146pi/512
   sin[147]  =  10'b1100110111;     //147pi/512
   cos[147]  =  10'b0010011110;     //147pi/512
   sin[148]  =  10'b1100110110;     //148pi/512
   cos[148]  =  10'b0010011101;     //148pi/512
   sin[149]  =  10'b1100110101;     //149pi/512
   cos[149]  =  10'b0010011100;     //149pi/512
   sin[150]  =  10'b1100110100;     //150pi/512
   cos[150]  =  10'b0010011011;     //150pi/512
   sin[151]  =  10'b1100110011;     //151pi/512
   cos[151]  =  10'b0010011001;     //151pi/512
   sin[152]  =  10'b1100110010;     //152pi/512
   cos[152]  =  10'b0010011000;     //152pi/512
   sin[153]  =  10'b1100110001;     //153pi/512
   cos[153]  =  10'b0010010111;     //153pi/512
   sin[154]  =  10'b1100110001;     //154pi/512
   cos[154]  =  10'b0010010101;     //154pi/512
   sin[155]  =  10'b1100110000;     //155pi/512
   cos[155]  =  10'b0010010100;     //155pi/512
   sin[156]  =  10'b1100101111;     //156pi/512
   cos[156]  =  10'b0010010011;     //156pi/512
   sin[157]  =  10'b1100101110;     //157pi/512
   cos[157]  =  10'b0010010010;     //157pi/512
   sin[158]  =  10'b1100101101;     //158pi/512
   cos[158]  =  10'b0010010000;     //158pi/512
   sin[159]  =  10'b1100101100;     //159pi/512
   cos[159]  =  10'b0010001111;     //159pi/512
   sin[160]  =  10'b1100101011;     //160pi/512
   cos[160]  =  10'b0010001110;     //160pi/512
   sin[161]  =  10'b1100101010;     //161pi/512
   cos[161]  =  10'b0010001100;     //161pi/512
   sin[162]  =  10'b1100101001;     //162pi/512
   cos[162]  =  10'b0010001011;     //162pi/512
   sin[163]  =  10'b1100101001;     //163pi/512
   cos[163]  =  10'b0010001010;     //163pi/512
   sin[164]  =  10'b1100101000;     //164pi/512
   cos[164]  =  10'b0010001000;     //164pi/512
   sin[165]  =  10'b1100100111;     //165pi/512
   cos[165]  =  10'b0010000111;     //165pi/512
   sin[166]  =  10'b1100100110;     //166pi/512
   cos[166]  =  10'b0010000110;     //166pi/512
   sin[167]  =  10'b1100100101;     //167pi/512
   cos[167]  =  10'b0010000100;     //167pi/512
   sin[168]  =  10'b1100100100;     //168pi/512
   cos[168]  =  10'b0010000011;     //168pi/512
   sin[169]  =  10'b1100100100;     //169pi/512
   cos[169]  =  10'b0010000010;     //169pi/512
   sin[170]  =  10'b1100100011;     //170pi/512
   cos[170]  =  10'b0010000000;     //170pi/512
   sin[171]  =  10'b1100100010;     //171pi/512
   cos[171]  =  10'b0001111111;     //171pi/512
   sin[172]  =  10'b1100100001;     //172pi/512
   cos[172]  =  10'b0001111110;     //172pi/512
   sin[173]  =  10'b1100100000;     //173pi/512
   cos[173]  =  10'b0001111100;     //173pi/512
   sin[174]  =  10'b1100100000;     //174pi/512
   cos[174]  =  10'b0001111011;     //174pi/512
   sin[175]  =  10'b1100011111;     //175pi/512
   cos[175]  =  10'b0001111010;     //175pi/512
   sin[176]  =  10'b1100011110;     //176pi/512
   cos[176]  =  10'b0001111000;     //176pi/512
   sin[177]  =  10'b1100011101;     //177pi/512
   cos[177]  =  10'b0001110111;     //177pi/512
   sin[178]  =  10'b1100011101;     //178pi/512
   cos[178]  =  10'b0001110101;     //178pi/512
   sin[179]  =  10'b1100011100;     //179pi/512
   cos[179]  =  10'b0001110100;     //179pi/512
   sin[180]  =  10'b1100011011;     //180pi/512
   cos[180]  =  10'b0001110011;     //180pi/512
   sin[181]  =  10'b1100011011;     //181pi/512
   cos[181]  =  10'b0001110001;     //181pi/512
   sin[182]  =  10'b1100011010;     //182pi/512
   cos[182]  =  10'b0001110000;     //182pi/512
   sin[183]  =  10'b1100011001;     //183pi/512
   cos[183]  =  10'b0001101110;     //183pi/512
   sin[184]  =  10'b1100011001;     //184pi/512
   cos[184]  =  10'b0001101101;     //184pi/512
   sin[185]  =  10'b1100011000;     //185pi/512
   cos[185]  =  10'b0001101100;     //185pi/512
   sin[186]  =  10'b1100010111;     //186pi/512
   cos[186]  =  10'b0001101010;     //186pi/512
   sin[187]  =  10'b1100010111;     //187pi/512
   cos[187]  =  10'b0001101001;     //187pi/512
   sin[188]  =  10'b1100010110;     //188pi/512
   cos[188]  =  10'b0001100111;     //188pi/512
   sin[189]  =  10'b1100010101;     //189pi/512
   cos[189]  =  10'b0001100110;     //189pi/512
   sin[190]  =  10'b1100010101;     //190pi/512
   cos[190]  =  10'b0001100100;     //190pi/512
   sin[191]  =  10'b1100010100;     //191pi/512
   cos[191]  =  10'b0001100011;     //191pi/512
   sin[192]  =  10'b1100010011;     //192pi/512
   cos[192]  =  10'b0001100001;     //192pi/512
   sin[193]  =  10'b1100010011;     //193pi/512
   cos[193]  =  10'b0001100000;     //193pi/512
   sin[194]  =  10'b1100010010;     //194pi/512
   cos[194]  =  10'b0001011111;     //194pi/512
   sin[195]  =  10'b1100010010;     //195pi/512
   cos[195]  =  10'b0001011101;     //195pi/512
   sin[196]  =  10'b1100010001;     //196pi/512
   cos[196]  =  10'b0001011100;     //196pi/512
   sin[197]  =  10'b1100010001;     //197pi/512
   cos[197]  =  10'b0001011010;     //197pi/512
   sin[198]  =  10'b1100010000;     //198pi/512
   cos[198]  =  10'b0001011001;     //198pi/512
   sin[199]  =  10'b1100001111;     //199pi/512
   cos[199]  =  10'b0001010111;     //199pi/512
   sin[200]  =  10'b1100001111;     //200pi/512
   cos[200]  =  10'b0001010110;     //200pi/512
   sin[201]  =  10'b1100001110;     //201pi/512
   cos[201]  =  10'b0001010100;     //201pi/512
   sin[202]  =  10'b1100001110;     //202pi/512
   cos[202]  =  10'b0001010011;     //202pi/512
   sin[203]  =  10'b1100001101;     //203pi/512
   cos[203]  =  10'b0001010001;     //203pi/512
   sin[204]  =  10'b1100001101;     //204pi/512
   cos[204]  =  10'b0001010000;     //204pi/512
   sin[205]  =  10'b1100001100;     //205pi/512
   cos[205]  =  10'b0001001110;     //205pi/512
   sin[206]  =  10'b1100001100;     //206pi/512
   cos[206]  =  10'b0001001101;     //206pi/512
   sin[207]  =  10'b1100001011;     //207pi/512
   cos[207]  =  10'b0001001011;     //207pi/512
   sin[208]  =  10'b1100001011;     //208pi/512
   cos[208]  =  10'b0001001010;     //208pi/512
   sin[209]  =  10'b1100001011;     //209pi/512
   cos[209]  =  10'b0001001000;     //209pi/512
   sin[210]  =  10'b1100001010;     //210pi/512
   cos[210]  =  10'b0001000111;     //210pi/512
   sin[211]  =  10'b1100001010;     //211pi/512
   cos[211]  =  10'b0001000101;     //211pi/512
   sin[212]  =  10'b1100001001;     //212pi/512
   cos[212]  =  10'b0001000100;     //212pi/512
   sin[213]  =  10'b1100001001;     //213pi/512
   cos[213]  =  10'b0001000010;     //213pi/512
   sin[214]  =  10'b1100001000;     //214pi/512
   cos[214]  =  10'b0001000001;     //214pi/512
   sin[215]  =  10'b1100001000;     //215pi/512
   cos[215]  =  10'b0000111111;     //215pi/512
   sin[216]  =  10'b1100001000;     //216pi/512
   cos[216]  =  10'b0000111110;     //216pi/512
   sin[217]  =  10'b1100000111;     //217pi/512
   cos[217]  =  10'b0000111100;     //217pi/512
   sin[218]  =  10'b1100000111;     //218pi/512
   cos[218]  =  10'b0000111011;     //218pi/512
   sin[219]  =  10'b1100000111;     //219pi/512
   cos[219]  =  10'b0000111001;     //219pi/512
   sin[220]  =  10'b1100000110;     //220pi/512
   cos[220]  =  10'b0000111000;     //220pi/512
   sin[221]  =  10'b1100000110;     //221pi/512
   cos[221]  =  10'b0000110110;     //221pi/512
   sin[222]  =  10'b1100000110;     //222pi/512
   cos[222]  =  10'b0000110101;     //222pi/512
   sin[223]  =  10'b1100000101;     //223pi/512
   cos[223]  =  10'b0000110011;     //223pi/512
   sin[224]  =  10'b1100000101;     //224pi/512
   cos[224]  =  10'b0000110001;     //224pi/512
   sin[225]  =  10'b1100000101;     //225pi/512
   cos[225]  =  10'b0000110000;     //225pi/512
   sin[226]  =  10'b1100000100;     //226pi/512
   cos[226]  =  10'b0000101110;     //226pi/512
   sin[227]  =  10'b1100000100;     //227pi/512
   cos[227]  =  10'b0000101101;     //227pi/512
   sin[228]  =  10'b1100000100;     //228pi/512
   cos[228]  =  10'b0000101011;     //228pi/512
   sin[229]  =  10'b1100000100;     //229pi/512
   cos[229]  =  10'b0000101010;     //229pi/512
   sin[230]  =  10'b1100000011;     //230pi/512
   cos[230]  =  10'b0000101000;     //230pi/512
   sin[231]  =  10'b1100000011;     //231pi/512
   cos[231]  =  10'b0000100111;     //231pi/512
   sin[232]  =  10'b1100000011;     //232pi/512
   cos[232]  =  10'b0000100101;     //232pi/512
   sin[233]  =  10'b1100000011;     //233pi/512
   cos[233]  =  10'b0000100100;     //233pi/512
   sin[234]  =  10'b1100000010;     //234pi/512
   cos[234]  =  10'b0000100010;     //234pi/512
   sin[235]  =  10'b1100000010;     //235pi/512
   cos[235]  =  10'b0000100000;     //235pi/512
   sin[236]  =  10'b1100000010;     //236pi/512
   cos[236]  =  10'b0000011111;     //236pi/512
   sin[237]  =  10'b1100000010;     //237pi/512
   cos[237]  =  10'b0000011101;     //237pi/512
   sin[238]  =  10'b1100000010;     //238pi/512
   cos[238]  =  10'b0000011100;     //238pi/512
   sin[239]  =  10'b1100000001;     //239pi/512
   cos[239]  =  10'b0000011010;     //239pi/512
   sin[240]  =  10'b1100000001;     //240pi/512
   cos[240]  =  10'b0000011001;     //240pi/512
   sin[241]  =  10'b1100000001;     //241pi/512
   cos[241]  =  10'b0000010111;     //241pi/512
   sin[242]  =  10'b1100000001;     //242pi/512
   cos[242]  =  10'b0000010101;     //242pi/512
   sin[243]  =  10'b1100000001;     //243pi/512
   cos[243]  =  10'b0000010100;     //243pi/512
   sin[244]  =  10'b1100000001;     //244pi/512
   cos[244]  =  10'b0000010010;     //244pi/512
   sin[245]  =  10'b1100000001;     //245pi/512
   cos[245]  =  10'b0000010001;     //245pi/512
   sin[246]  =  10'b1100000000;     //246pi/512
   cos[246]  =  10'b0000001111;     //246pi/512
   sin[247]  =  10'b1100000000;     //247pi/512
   cos[247]  =  10'b0000001110;     //247pi/512
   sin[248]  =  10'b1100000000;     //248pi/512
   cos[248]  =  10'b0000001100;     //248pi/512
   sin[249]  =  10'b1100000000;     //249pi/512
   cos[249]  =  10'b0000001010;     //249pi/512
   sin[250]  =  10'b1100000000;     //250pi/512
   cos[250]  =  10'b0000001001;     //250pi/512
   sin[251]  =  10'b1100000000;     //251pi/512
   cos[251]  =  10'b0000000111;     //251pi/512
   sin[252]  =  10'b1100000000;     //252pi/512
   cos[252]  =  10'b0000000110;     //252pi/512
   sin[253]  =  10'b1100000000;     //253pi/512
   cos[253]  =  10'b0000000100;     //253pi/512
   sin[254]  =  10'b1100000000;     //254pi/512
   cos[254]  =  10'b0000000011;     //254pi/512
   sin[255]  =  10'b1100000000;     //255pi/512
   cos[255]  =  10'b0000000001;     //255pi/512
   sin[256]  =  10'b1100000000;     //256pi/512
   cos[256]  =  10'b0000000000;     //256pi/512
   sin[257]  =  10'b1100000000;     //257pi/512
   cos[257]  =  10'b1111111110;     //257pi/512
   sin[258]  =  10'b1100000000;     //258pi/512
   cos[258]  =  10'b1111111101;     //258pi/512
   sin[259]  =  10'b1100000000;     //259pi/512
   cos[259]  =  10'b1111111011;     //259pi/512
   sin[260]  =  10'b1100000000;     //260pi/512
   cos[260]  =  10'b1111111010;     //260pi/512
   sin[261]  =  10'b1100000000;     //261pi/512
   cos[261]  =  10'b1111111000;     //261pi/512
   sin[262]  =  10'b1100000000;     //262pi/512
   cos[262]  =  10'b1111110111;     //262pi/512
   sin[263]  =  10'b1100000000;     //263pi/512
   cos[263]  =  10'b1111110101;     //263pi/512
   sin[264]  =  10'b1100000000;     //264pi/512
   cos[264]  =  10'b1111110011;     //264pi/512
   sin[265]  =  10'b1100000000;     //265pi/512
   cos[265]  =  10'b1111110010;     //265pi/512
   sin[266]  =  10'b1100000000;     //266pi/512
   cos[266]  =  10'b1111110000;     //266pi/512
   sin[267]  =  10'b1100000001;     //267pi/512
   cos[267]  =  10'b1111101111;     //267pi/512
   sin[268]  =  10'b1100000001;     //268pi/512
   cos[268]  =  10'b1111101101;     //268pi/512
   sin[269]  =  10'b1100000001;     //269pi/512
   cos[269]  =  10'b1111101100;     //269pi/512
   sin[270]  =  10'b1100000001;     //270pi/512
   cos[270]  =  10'b1111101010;     //270pi/512
   sin[271]  =  10'b1100000001;     //271pi/512
   cos[271]  =  10'b1111101000;     //271pi/512
   sin[272]  =  10'b1100000001;     //272pi/512
   cos[272]  =  10'b1111100111;     //272pi/512
   sin[273]  =  10'b1100000001;     //273pi/512
   cos[273]  =  10'b1111100101;     //273pi/512
   sin[274]  =  10'b1100000010;     //274pi/512
   cos[274]  =  10'b1111100100;     //274pi/512
   sin[275]  =  10'b1100000010;     //275pi/512
   cos[275]  =  10'b1111100010;     //275pi/512
   sin[276]  =  10'b1100000010;     //276pi/512
   cos[276]  =  10'b1111100001;     //276pi/512
   sin[277]  =  10'b1100000010;     //277pi/512
   cos[277]  =  10'b1111011111;     //277pi/512
   sin[278]  =  10'b1100000010;     //278pi/512
   cos[278]  =  10'b1111011110;     //278pi/512
   sin[279]  =  10'b1100000011;     //279pi/512
   cos[279]  =  10'b1111011100;     //279pi/512
   sin[280]  =  10'b1100000011;     //280pi/512
   cos[280]  =  10'b1111011010;     //280pi/512
   sin[281]  =  10'b1100000011;     //281pi/512
   cos[281]  =  10'b1111011001;     //281pi/512
   sin[282]  =  10'b1100000011;     //282pi/512
   cos[282]  =  10'b1111010111;     //282pi/512
   sin[283]  =  10'b1100000100;     //283pi/512
   cos[283]  =  10'b1111010110;     //283pi/512
   sin[284]  =  10'b1100000100;     //284pi/512
   cos[284]  =  10'b1111010100;     //284pi/512
   sin[285]  =  10'b1100000100;     //285pi/512
   cos[285]  =  10'b1111010011;     //285pi/512
   sin[286]  =  10'b1100000100;     //286pi/512
   cos[286]  =  10'b1111010001;     //286pi/512
   sin[287]  =  10'b1100000101;     //287pi/512
   cos[287]  =  10'b1111010000;     //287pi/512
   sin[288]  =  10'b1100000101;     //288pi/512
   cos[288]  =  10'b1111001110;     //288pi/512
   sin[289]  =  10'b1100000101;     //289pi/512
   cos[289]  =  10'b1111001101;     //289pi/512
   sin[290]  =  10'b1100000110;     //290pi/512
   cos[290]  =  10'b1111001011;     //290pi/512
   sin[291]  =  10'b1100000110;     //291pi/512
   cos[291]  =  10'b1111001001;     //291pi/512
   sin[292]  =  10'b1100000110;     //292pi/512
   cos[292]  =  10'b1111001000;     //292pi/512
   sin[293]  =  10'b1100000111;     //293pi/512
   cos[293]  =  10'b1111000110;     //293pi/512
   sin[294]  =  10'b1100000111;     //294pi/512
   cos[294]  =  10'b1111000101;     //294pi/512
   sin[295]  =  10'b1100000111;     //295pi/512
   cos[295]  =  10'b1111000011;     //295pi/512
   sin[296]  =  10'b1100001000;     //296pi/512
   cos[296]  =  10'b1111000010;     //296pi/512
   sin[297]  =  10'b1100001000;     //297pi/512
   cos[297]  =  10'b1111000000;     //297pi/512
   sin[298]  =  10'b1100001000;     //298pi/512
   cos[298]  =  10'b1110111111;     //298pi/512
   sin[299]  =  10'b1100001001;     //299pi/512
   cos[299]  =  10'b1110111101;     //299pi/512
   sin[300]  =  10'b1100001001;     //300pi/512
   cos[300]  =  10'b1110111100;     //300pi/512
   sin[301]  =  10'b1100001010;     //301pi/512
   cos[301]  =  10'b1110111010;     //301pi/512
   sin[302]  =  10'b1100001010;     //302pi/512
   cos[302]  =  10'b1110111001;     //302pi/512
   sin[303]  =  10'b1100001011;     //303pi/512
   cos[303]  =  10'b1110110111;     //303pi/512
   sin[304]  =  10'b1100001011;     //304pi/512
   cos[304]  =  10'b1110110110;     //304pi/512
   sin[305]  =  10'b1100001011;     //305pi/512
   cos[305]  =  10'b1110110100;     //305pi/512
   sin[306]  =  10'b1100001100;     //306pi/512
   cos[306]  =  10'b1110110011;     //306pi/512
   sin[307]  =  10'b1100001100;     //307pi/512
   cos[307]  =  10'b1110110001;     //307pi/512
   sin[308]  =  10'b1100001101;     //308pi/512
   cos[308]  =  10'b1110110000;     //308pi/512
   sin[309]  =  10'b1100001101;     //309pi/512
   cos[309]  =  10'b1110101110;     //309pi/512
   sin[310]  =  10'b1100001110;     //310pi/512
   cos[310]  =  10'b1110101101;     //310pi/512
   sin[311]  =  10'b1100001110;     //311pi/512
   cos[311]  =  10'b1110101011;     //311pi/512
   sin[312]  =  10'b1100001111;     //312pi/512
   cos[312]  =  10'b1110101010;     //312pi/512
   sin[313]  =  10'b1100001111;     //313pi/512
   cos[313]  =  10'b1110101000;     //313pi/512
   sin[314]  =  10'b1100010000;     //314pi/512
   cos[314]  =  10'b1110100111;     //314pi/512
   sin[315]  =  10'b1100010001;     //315pi/512
   cos[315]  =  10'b1110100101;     //315pi/512
   sin[316]  =  10'b1100010001;     //316pi/512
   cos[316]  =  10'b1110100100;     //316pi/512
   sin[317]  =  10'b1100010010;     //317pi/512
   cos[317]  =  10'b1110100010;     //317pi/512
   sin[318]  =  10'b1100010010;     //318pi/512
   cos[318]  =  10'b1110100001;     //318pi/512
   sin[319]  =  10'b1100010011;     //319pi/512
   cos[319]  =  10'b1110011111;     //319pi/512
   sin[320]  =  10'b1100010011;     //320pi/512
   cos[320]  =  10'b1110011110;     //320pi/512
   sin[321]  =  10'b1100010100;     //321pi/512
   cos[321]  =  10'b1110011101;     //321pi/512
   sin[322]  =  10'b1100010101;     //322pi/512
   cos[322]  =  10'b1110011011;     //322pi/512
   sin[323]  =  10'b1100010101;     //323pi/512
   cos[323]  =  10'b1110011010;     //323pi/512
   sin[324]  =  10'b1100010110;     //324pi/512
   cos[324]  =  10'b1110011000;     //324pi/512
   sin[325]  =  10'b1100010111;     //325pi/512
   cos[325]  =  10'b1110010111;     //325pi/512
   sin[326]  =  10'b1100010111;     //326pi/512
   cos[326]  =  10'b1110010101;     //326pi/512
   sin[327]  =  10'b1100011000;     //327pi/512
   cos[327]  =  10'b1110010100;     //327pi/512
   sin[328]  =  10'b1100011001;     //328pi/512
   cos[328]  =  10'b1110010011;     //328pi/512
   sin[329]  =  10'b1100011001;     //329pi/512
   cos[329]  =  10'b1110010001;     //329pi/512
   sin[330]  =  10'b1100011010;     //330pi/512
   cos[330]  =  10'b1110010000;     //330pi/512
   sin[331]  =  10'b1100011011;     //331pi/512
   cos[331]  =  10'b1110001110;     //331pi/512
   sin[332]  =  10'b1100011011;     //332pi/512
   cos[332]  =  10'b1110001101;     //332pi/512
   sin[333]  =  10'b1100011100;     //333pi/512
   cos[333]  =  10'b1110001011;     //333pi/512
   sin[334]  =  10'b1100011101;     //334pi/512
   cos[334]  =  10'b1110001010;     //334pi/512
   sin[335]  =  10'b1100011101;     //335pi/512
   cos[335]  =  10'b1110001001;     //335pi/512
   sin[336]  =  10'b1100011110;     //336pi/512
   cos[336]  =  10'b1110000111;     //336pi/512
   sin[337]  =  10'b1100011111;     //337pi/512
   cos[337]  =  10'b1110000110;     //337pi/512
   sin[338]  =  10'b1100100000;     //338pi/512
   cos[338]  =  10'b1110000101;     //338pi/512
   sin[339]  =  10'b1100100000;     //339pi/512
   cos[339]  =  10'b1110000011;     //339pi/512
   sin[340]  =  10'b1100100001;     //340pi/512
   cos[340]  =  10'b1110000010;     //340pi/512
   sin[341]  =  10'b1100100010;     //341pi/512
   cos[341]  =  10'b1110000000;     //341pi/512
   sin[342]  =  10'b1100100011;     //342pi/512
   cos[342]  =  10'b1101111111;     //342pi/512
   sin[343]  =  10'b1100100100;     //343pi/512
   cos[343]  =  10'b1101111110;     //343pi/512
   sin[344]  =  10'b1100100100;     //344pi/512
   cos[344]  =  10'b1101111100;     //344pi/512
   sin[345]  =  10'b1100100101;     //345pi/512
   cos[345]  =  10'b1101111011;     //345pi/512
   sin[346]  =  10'b1100100110;     //346pi/512
   cos[346]  =  10'b1101111010;     //346pi/512
   sin[347]  =  10'b1100100111;     //347pi/512
   cos[347]  =  10'b1101111000;     //347pi/512
   sin[348]  =  10'b1100101000;     //348pi/512
   cos[348]  =  10'b1101110111;     //348pi/512
   sin[349]  =  10'b1100101001;     //349pi/512
   cos[349]  =  10'b1101110110;     //349pi/512
   sin[350]  =  10'b1100101001;     //350pi/512
   cos[350]  =  10'b1101110100;     //350pi/512
   sin[351]  =  10'b1100101010;     //351pi/512
   cos[351]  =  10'b1101110011;     //351pi/512
   sin[352]  =  10'b1100101011;     //352pi/512
   cos[352]  =  10'b1101110010;     //352pi/512
   sin[353]  =  10'b1100101100;     //353pi/512
   cos[353]  =  10'b1101110000;     //353pi/512
   sin[354]  =  10'b1100101101;     //354pi/512
   cos[354]  =  10'b1101101111;     //354pi/512
   sin[355]  =  10'b1100101110;     //355pi/512
   cos[355]  =  10'b1101101110;     //355pi/512
   sin[356]  =  10'b1100101111;     //356pi/512
   cos[356]  =  10'b1101101101;     //356pi/512
   sin[357]  =  10'b1100110000;     //357pi/512
   cos[357]  =  10'b1101101011;     //357pi/512
   sin[358]  =  10'b1100110001;     //358pi/512
   cos[358]  =  10'b1101101010;     //358pi/512
   sin[359]  =  10'b1100110001;     //359pi/512
   cos[359]  =  10'b1101101001;     //359pi/512
   sin[360]  =  10'b1100110010;     //360pi/512
   cos[360]  =  10'b1101101000;     //360pi/512
   sin[361]  =  10'b1100110011;     //361pi/512
   cos[361]  =  10'b1101100110;     //361pi/512
   sin[362]  =  10'b1100110100;     //362pi/512
   cos[362]  =  10'b1101100101;     //362pi/512
   sin[363]  =  10'b1100110101;     //363pi/512
   cos[363]  =  10'b1101100100;     //363pi/512
   sin[364]  =  10'b1100110110;     //364pi/512
   cos[364]  =  10'b1101100011;     //364pi/512
   sin[365]  =  10'b1100110111;     //365pi/512
   cos[365]  =  10'b1101100001;     //365pi/512
   sin[366]  =  10'b1100111000;     //366pi/512
   cos[366]  =  10'b1101100000;     //366pi/512
   sin[367]  =  10'b1100111001;     //367pi/512
   cos[367]  =  10'b1101011111;     //367pi/512
   sin[368]  =  10'b1100111010;     //368pi/512
   cos[368]  =  10'b1101011110;     //368pi/512
   sin[369]  =  10'b1100111011;     //369pi/512
   cos[369]  =  10'b1101011100;     //369pi/512
   sin[370]  =  10'b1100111100;     //370pi/512
   cos[370]  =  10'b1101011011;     //370pi/512
   sin[371]  =  10'b1100111101;     //371pi/512
   cos[371]  =  10'b1101011010;     //371pi/512
   sin[372]  =  10'b1100111110;     //372pi/512
   cos[372]  =  10'b1101011001;     //372pi/512
   sin[373]  =  10'b1100111111;     //373pi/512
   cos[373]  =  10'b1101011000;     //373pi/512
   sin[374]  =  10'b1101000000;     //374pi/512
   cos[374]  =  10'b1101010110;     //374pi/512
   sin[375]  =  10'b1101000001;     //375pi/512
   cos[375]  =  10'b1101010101;     //375pi/512
   sin[376]  =  10'b1101000010;     //376pi/512
   cos[376]  =  10'b1101010100;     //376pi/512
   sin[377]  =  10'b1101000011;     //377pi/512
   cos[377]  =  10'b1101010011;     //377pi/512
   sin[378]  =  10'b1101000100;     //378pi/512
   cos[378]  =  10'b1101010010;     //378pi/512
   sin[379]  =  10'b1101000110;     //379pi/512
   cos[379]  =  10'b1101010001;     //379pi/512
   sin[380]  =  10'b1101000111;     //380pi/512
   cos[380]  =  10'b1101001111;     //380pi/512
   sin[381]  =  10'b1101001000;     //381pi/512
   cos[381]  =  10'b1101001110;     //381pi/512
   sin[382]  =  10'b1101001001;     //382pi/512
   cos[382]  =  10'b1101001101;     //382pi/512
   sin[383]  =  10'b1101001010;     //383pi/512
   cos[383]  =  10'b1101001100;     //383pi/512
   sin[384]  =  10'b1101001011;     //384pi/512
   cos[384]  =  10'b1101001011;     //384pi/512
   sin[385]  =  10'b1101001100;     //385pi/512
   cos[385]  =  10'b1101001010;     //385pi/512
   sin[386]  =  10'b1101001101;     //386pi/512
   cos[386]  =  10'b1101001001;     //386pi/512
   sin[387]  =  10'b1101001110;     //387pi/512
   cos[387]  =  10'b1101001000;     //387pi/512
   sin[388]  =  10'b1101001111;     //388pi/512
   cos[388]  =  10'b1101000111;     //388pi/512
   sin[389]  =  10'b1101010001;     //389pi/512
   cos[389]  =  10'b1101000110;     //389pi/512
   sin[390]  =  10'b1101010010;     //390pi/512
   cos[390]  =  10'b1101000100;     //390pi/512
   sin[391]  =  10'b1101010011;     //391pi/512
   cos[391]  =  10'b1101000011;     //391pi/512
   sin[392]  =  10'b1101010100;     //392pi/512
   cos[392]  =  10'b1101000010;     //392pi/512
   sin[393]  =  10'b1101010101;     //393pi/512
   cos[393]  =  10'b1101000001;     //393pi/512
   sin[394]  =  10'b1101010110;     //394pi/512
   cos[394]  =  10'b1101000000;     //394pi/512
   sin[395]  =  10'b1101011000;     //395pi/512
   cos[395]  =  10'b1100111111;     //395pi/512
   sin[396]  =  10'b1101011001;     //396pi/512
   cos[396]  =  10'b1100111110;     //396pi/512
   sin[397]  =  10'b1101011010;     //397pi/512
   cos[397]  =  10'b1100111101;     //397pi/512
   sin[398]  =  10'b1101011011;     //398pi/512
   cos[398]  =  10'b1100111100;     //398pi/512
   sin[399]  =  10'b1101011100;     //399pi/512
   cos[399]  =  10'b1100111011;     //399pi/512
   sin[400]  =  10'b1101011110;     //400pi/512
   cos[400]  =  10'b1100111010;     //400pi/512
   sin[401]  =  10'b1101011111;     //401pi/512
   cos[401]  =  10'b1100111001;     //401pi/512
   sin[402]  =  10'b1101100000;     //402pi/512
   cos[402]  =  10'b1100111000;     //402pi/512
   sin[403]  =  10'b1101100001;     //403pi/512
   cos[403]  =  10'b1100110111;     //403pi/512
   sin[404]  =  10'b1101100011;     //404pi/512
   cos[404]  =  10'b1100110110;     //404pi/512
   sin[405]  =  10'b1101100100;     //405pi/512
   cos[405]  =  10'b1100110101;     //405pi/512
   sin[406]  =  10'b1101100101;     //406pi/512
   cos[406]  =  10'b1100110100;     //406pi/512
   sin[407]  =  10'b1101100110;     //407pi/512
   cos[407]  =  10'b1100110011;     //407pi/512
   sin[408]  =  10'b1101101000;     //408pi/512
   cos[408]  =  10'b1100110010;     //408pi/512
   sin[409]  =  10'b1101101001;     //409pi/512
   cos[409]  =  10'b1100110001;     //409pi/512
   sin[410]  =  10'b1101101010;     //410pi/512
   cos[410]  =  10'b1100110001;     //410pi/512
   sin[411]  =  10'b1101101011;     //411pi/512
   cos[411]  =  10'b1100110000;     //411pi/512
   sin[412]  =  10'b1101101101;     //412pi/512
   cos[412]  =  10'b1100101111;     //412pi/512
   sin[413]  =  10'b1101101110;     //413pi/512
   cos[413]  =  10'b1100101110;     //413pi/512
   sin[414]  =  10'b1101101111;     //414pi/512
   cos[414]  =  10'b1100101101;     //414pi/512
   sin[415]  =  10'b1101110000;     //415pi/512
   cos[415]  =  10'b1100101100;     //415pi/512
   sin[416]  =  10'b1101110010;     //416pi/512
   cos[416]  =  10'b1100101011;     //416pi/512
   sin[417]  =  10'b1101110011;     //417pi/512
   cos[417]  =  10'b1100101010;     //417pi/512
   sin[418]  =  10'b1101110100;     //418pi/512
   cos[418]  =  10'b1100101001;     //418pi/512
   sin[419]  =  10'b1101110110;     //419pi/512
   cos[419]  =  10'b1100101001;     //419pi/512
   sin[420]  =  10'b1101110111;     //420pi/512
   cos[420]  =  10'b1100101000;     //420pi/512
   sin[421]  =  10'b1101111000;     //421pi/512
   cos[421]  =  10'b1100100111;     //421pi/512
   sin[422]  =  10'b1101111010;     //422pi/512
   cos[422]  =  10'b1100100110;     //422pi/512
   sin[423]  =  10'b1101111011;     //423pi/512
   cos[423]  =  10'b1100100101;     //423pi/512
   sin[424]  =  10'b1101111100;     //424pi/512
   cos[424]  =  10'b1100100100;     //424pi/512
   sin[425]  =  10'b1101111110;     //425pi/512
   cos[425]  =  10'b1100100100;     //425pi/512
   sin[426]  =  10'b1101111111;     //426pi/512
   cos[426]  =  10'b1100100011;     //426pi/512
   sin[427]  =  10'b1110000000;     //427pi/512
   cos[427]  =  10'b1100100010;     //427pi/512
   sin[428]  =  10'b1110000010;     //428pi/512
   cos[428]  =  10'b1100100001;     //428pi/512
   sin[429]  =  10'b1110000011;     //429pi/512
   cos[429]  =  10'b1100100000;     //429pi/512
   sin[430]  =  10'b1110000101;     //430pi/512
   cos[430]  =  10'b1100100000;     //430pi/512
   sin[431]  =  10'b1110000110;     //431pi/512
   cos[431]  =  10'b1100011111;     //431pi/512
   sin[432]  =  10'b1110000111;     //432pi/512
   cos[432]  =  10'b1100011110;     //432pi/512
   sin[433]  =  10'b1110001001;     //433pi/512
   cos[433]  =  10'b1100011101;     //433pi/512
   sin[434]  =  10'b1110001010;     //434pi/512
   cos[434]  =  10'b1100011101;     //434pi/512
   sin[435]  =  10'b1110001011;     //435pi/512
   cos[435]  =  10'b1100011100;     //435pi/512
   sin[436]  =  10'b1110001101;     //436pi/512
   cos[436]  =  10'b1100011011;     //436pi/512
   sin[437]  =  10'b1110001110;     //437pi/512
   cos[437]  =  10'b1100011011;     //437pi/512
   sin[438]  =  10'b1110010000;     //438pi/512
   cos[438]  =  10'b1100011010;     //438pi/512
   sin[439]  =  10'b1110010001;     //439pi/512
   cos[439]  =  10'b1100011001;     //439pi/512
   sin[440]  =  10'b1110010011;     //440pi/512
   cos[440]  =  10'b1100011001;     //440pi/512
   sin[441]  =  10'b1110010100;     //441pi/512
   cos[441]  =  10'b1100011000;     //441pi/512
   sin[442]  =  10'b1110010101;     //442pi/512
   cos[442]  =  10'b1100010111;     //442pi/512
   sin[443]  =  10'b1110010111;     //443pi/512
   cos[443]  =  10'b1100010111;     //443pi/512
   sin[444]  =  10'b1110011000;     //444pi/512
   cos[444]  =  10'b1100010110;     //444pi/512
   sin[445]  =  10'b1110011010;     //445pi/512
   cos[445]  =  10'b1100010101;     //445pi/512
   sin[446]  =  10'b1110011011;     //446pi/512
   cos[446]  =  10'b1100010101;     //446pi/512
   sin[447]  =  10'b1110011101;     //447pi/512
   cos[447]  =  10'b1100010100;     //447pi/512
   sin[448]  =  10'b1110011110;     //448pi/512
   cos[448]  =  10'b1100010011;     //448pi/512
   sin[449]  =  10'b1110011111;     //449pi/512
   cos[449]  =  10'b1100010011;     //449pi/512
   sin[450]  =  10'b1110100001;     //450pi/512
   cos[450]  =  10'b1100010010;     //450pi/512
   sin[451]  =  10'b1110100010;     //451pi/512
   cos[451]  =  10'b1100010010;     //451pi/512
   sin[452]  =  10'b1110100100;     //452pi/512
   cos[452]  =  10'b1100010001;     //452pi/512
   sin[453]  =  10'b1110100101;     //453pi/512
   cos[453]  =  10'b1100010001;     //453pi/512
   sin[454]  =  10'b1110100111;     //454pi/512
   cos[454]  =  10'b1100010000;     //454pi/512
   sin[455]  =  10'b1110101000;     //455pi/512
   cos[455]  =  10'b1100001111;     //455pi/512
   sin[456]  =  10'b1110101010;     //456pi/512
   cos[456]  =  10'b1100001111;     //456pi/512
   sin[457]  =  10'b1110101011;     //457pi/512
   cos[457]  =  10'b1100001110;     //457pi/512
   sin[458]  =  10'b1110101101;     //458pi/512
   cos[458]  =  10'b1100001110;     //458pi/512
   sin[459]  =  10'b1110101110;     //459pi/512
   cos[459]  =  10'b1100001101;     //459pi/512
   sin[460]  =  10'b1110110000;     //460pi/512
   cos[460]  =  10'b1100001101;     //460pi/512
   sin[461]  =  10'b1110110001;     //461pi/512
   cos[461]  =  10'b1100001100;     //461pi/512
   sin[462]  =  10'b1110110011;     //462pi/512
   cos[462]  =  10'b1100001100;     //462pi/512
   sin[463]  =  10'b1110110100;     //463pi/512
   cos[463]  =  10'b1100001011;     //463pi/512
   sin[464]  =  10'b1110110110;     //464pi/512
   cos[464]  =  10'b1100001011;     //464pi/512
   sin[465]  =  10'b1110110111;     //465pi/512
   cos[465]  =  10'b1100001011;     //465pi/512
   sin[466]  =  10'b1110111001;     //466pi/512
   cos[466]  =  10'b1100001010;     //466pi/512
   sin[467]  =  10'b1110111010;     //467pi/512
   cos[467]  =  10'b1100001010;     //467pi/512
   sin[468]  =  10'b1110111100;     //468pi/512
   cos[468]  =  10'b1100001001;     //468pi/512
   sin[469]  =  10'b1110111101;     //469pi/512
   cos[469]  =  10'b1100001001;     //469pi/512
   sin[470]  =  10'b1110111111;     //470pi/512
   cos[470]  =  10'b1100001000;     //470pi/512
   sin[471]  =  10'b1111000000;     //471pi/512
   cos[471]  =  10'b1100001000;     //471pi/512
   sin[472]  =  10'b1111000010;     //472pi/512
   cos[472]  =  10'b1100001000;     //472pi/512
   sin[473]  =  10'b1111000011;     //473pi/512
   cos[473]  =  10'b1100000111;     //473pi/512
   sin[474]  =  10'b1111000101;     //474pi/512
   cos[474]  =  10'b1100000111;     //474pi/512
   sin[475]  =  10'b1111000110;     //475pi/512
   cos[475]  =  10'b1100000111;     //475pi/512
   sin[476]  =  10'b1111001000;     //476pi/512
   cos[476]  =  10'b1100000110;     //476pi/512
   sin[477]  =  10'b1111001001;     //477pi/512
   cos[477]  =  10'b1100000110;     //477pi/512
   sin[478]  =  10'b1111001011;     //478pi/512
   cos[478]  =  10'b1100000110;     //478pi/512
   sin[479]  =  10'b1111001101;     //479pi/512
   cos[479]  =  10'b1100000101;     //479pi/512
   sin[480]  =  10'b1111001110;     //480pi/512
   cos[480]  =  10'b1100000101;     //480pi/512
   sin[481]  =  10'b1111010000;     //481pi/512
   cos[481]  =  10'b1100000101;     //481pi/512
   sin[482]  =  10'b1111010001;     //482pi/512
   cos[482]  =  10'b1100000100;     //482pi/512
   sin[483]  =  10'b1111010011;     //483pi/512
   cos[483]  =  10'b1100000100;     //483pi/512
   sin[484]  =  10'b1111010100;     //484pi/512
   cos[484]  =  10'b1100000100;     //484pi/512
   sin[485]  =  10'b1111010110;     //485pi/512
   cos[485]  =  10'b1100000100;     //485pi/512
   sin[486]  =  10'b1111010111;     //486pi/512
   cos[486]  =  10'b1100000011;     //486pi/512
   sin[487]  =  10'b1111011001;     //487pi/512
   cos[487]  =  10'b1100000011;     //487pi/512
   sin[488]  =  10'b1111011010;     //488pi/512
   cos[488]  =  10'b1100000011;     //488pi/512
   sin[489]  =  10'b1111011100;     //489pi/512
   cos[489]  =  10'b1100000011;     //489pi/512
   sin[490]  =  10'b1111011110;     //490pi/512
   cos[490]  =  10'b1100000010;     //490pi/512
   sin[491]  =  10'b1111011111;     //491pi/512
   cos[491]  =  10'b1100000010;     //491pi/512
   sin[492]  =  10'b1111100001;     //492pi/512
   cos[492]  =  10'b1100000010;     //492pi/512
   sin[493]  =  10'b1111100010;     //493pi/512
   cos[493]  =  10'b1100000010;     //493pi/512
   sin[494]  =  10'b1111100100;     //494pi/512
   cos[494]  =  10'b1100000010;     //494pi/512
   sin[495]  =  10'b1111100101;     //495pi/512
   cos[495]  =  10'b1100000001;     //495pi/512
   sin[496]  =  10'b1111100111;     //496pi/512
   cos[496]  =  10'b1100000001;     //496pi/512
   sin[497]  =  10'b1111101000;     //497pi/512
   cos[497]  =  10'b1100000001;     //497pi/512
   sin[498]  =  10'b1111101010;     //498pi/512
   cos[498]  =  10'b1100000001;     //498pi/512
   sin[499]  =  10'b1111101100;     //499pi/512
   cos[499]  =  10'b1100000001;     //499pi/512
   sin[500]  =  10'b1111101101;     //500pi/512
   cos[500]  =  10'b1100000001;     //500pi/512
   sin[501]  =  10'b1111101111;     //501pi/512
   cos[501]  =  10'b1100000001;     //501pi/512
   sin[502]  =  10'b1111110000;     //502pi/512
   cos[502]  =  10'b1100000000;     //502pi/512
   sin[503]  =  10'b1111110010;     //503pi/512
   cos[503]  =  10'b1100000000;     //503pi/512
   sin[504]  =  10'b1111110011;     //504pi/512
   cos[504]  =  10'b1100000000;     //504pi/512
   sin[505]  =  10'b1111110101;     //505pi/512
   cos[505]  =  10'b1100000000;     //505pi/512
   sin[506]  =  10'b1111110111;     //506pi/512
   cos[506]  =  10'b1100000000;     //506pi/512
   sin[507]  =  10'b1111111000;     //507pi/512
   cos[507]  =  10'b1100000000;     //507pi/512
   sin[508]  =  10'b1111111010;     //508pi/512
   cos[508]  =  10'b1100000000;     //508pi/512
   sin[509]  =  10'b1111111011;     //509pi/512
   cos[509]  =  10'b1100000000;     //509pi/512
   sin[510]  =  10'b1111111101;     //510pi/512
   cos[510]  =  10'b1100000000;     //510pi/512
   sin[511]  =  10'b1111111110;     //511pi/512
   cos[511]  =  10'b1100000000;     //511pi/512

/////////////////////////////////////////////////////////////////

   m_sin[0]  =  10'b0000000000;     //0pi/512
   m_cos[0]  =  10'b0100000000;     //0pi/512
   m_sin[1]  =  10'b1111111111;     //1pi/512
   m_cos[1]  =  10'b0011111111;     //1pi/512
   m_sin[2]  =  10'b1111111101;     //2pi/512
   m_cos[2]  =  10'b0011111111;     //2pi/512
   m_sin[3]  =  10'b1111111100;     //3pi/512
   m_cos[3]  =  10'b0011111111;     //3pi/512
   m_sin[4]  =  10'b1111111011;     //4pi/512
   m_cos[4]  =  10'b0011111111;     //4pi/512
   m_sin[5]  =  10'b1111111010;     //5pi/512
   m_cos[5]  =  10'b0011111111;     //5pi/512
   m_sin[6]  =  10'b1111111000;     //6pi/512
   m_cos[6]  =  10'b0011111111;     //6pi/512
   m_sin[7]  =  10'b1111110111;     //7pi/512
   m_cos[7]  =  10'b0011111111;     //7pi/512
   m_sin[8]  =  10'b1111110110;     //8pi/512
   m_cos[8]  =  10'b0011111111;     //8pi/512
   m_sin[9]  =  10'b1111110101;     //9pi/512
   m_cos[9]  =  10'b0011111111;     //9pi/512
   m_sin[10]  =  10'b1111110011;     //10pi/512
   m_cos[10]  =  10'b0011111111;     //10pi/512
   m_sin[11]  =  10'b1111110010;     //11pi/512
   m_cos[11]  =  10'b0011111111;     //11pi/512
   m_sin[12]  =  10'b1111110001;     //12pi/512
   m_cos[12]  =  10'b0011111111;     //12pi/512
   m_sin[13]  =  10'b1111110000;     //13pi/512
   m_cos[13]  =  10'b0011111111;     //13pi/512
   m_sin[14]  =  10'b1111101110;     //14pi/512
   m_cos[14]  =  10'b0011111111;     //14pi/512
   m_sin[15]  =  10'b1111101101;     //15pi/512
   m_cos[15]  =  10'b0011111111;     //15pi/512
   m_sin[16]  =  10'b1111101100;     //16pi/512
   m_cos[16]  =  10'b0011111111;     //16pi/512
   m_sin[17]  =  10'b1111101011;     //17pi/512
   m_cos[17]  =  10'b0011111111;     //17pi/512
   m_sin[18]  =  10'b1111101001;     //18pi/512
   m_cos[18]  =  10'b0011111111;     //18pi/512
   m_sin[19]  =  10'b1111101000;     //19pi/512
   m_cos[19]  =  10'b0011111110;     //19pi/512
   m_sin[20]  =  10'b1111100111;     //20pi/512
   m_cos[20]  =  10'b0011111110;     //20pi/512
   m_sin[21]  =  10'b1111100110;     //21pi/512
   m_cos[21]  =  10'b0011111110;     //21pi/512
   m_sin[22]  =  10'b1111100100;     //22pi/512
   m_cos[22]  =  10'b0011111110;     //22pi/512
   m_sin[23]  =  10'b1111100011;     //23pi/512
   m_cos[23]  =  10'b0011111110;     //23pi/512
   m_sin[24]  =  10'b1111100010;     //24pi/512
   m_cos[24]  =  10'b0011111110;     //24pi/512
   m_sin[25]  =  10'b1111100001;     //25pi/512
   m_cos[25]  =  10'b0011111110;     //25pi/512
   m_sin[26]  =  10'b1111011111;     //26pi/512
   m_cos[26]  =  10'b0011111101;     //26pi/512
   m_sin[27]  =  10'b1111011110;     //27pi/512
   m_cos[27]  =  10'b0011111101;     //27pi/512
   m_sin[28]  =  10'b1111011101;     //28pi/512
   m_cos[28]  =  10'b0011111101;     //28pi/512
   m_sin[29]  =  10'b1111011100;     //29pi/512
   m_cos[29]  =  10'b0011111101;     //29pi/512
   m_sin[30]  =  10'b1111011010;     //30pi/512
   m_cos[30]  =  10'b0011111101;     //30pi/512
   m_sin[31]  =  10'b1111011001;     //31pi/512
   m_cos[31]  =  10'b0011111101;     //31pi/512
   m_sin[32]  =  10'b1111011000;     //32pi/512
   m_cos[32]  =  10'b0011111100;     //32pi/512
   m_sin[33]  =  10'b1111010111;     //33pi/512
   m_cos[33]  =  10'b0011111100;     //33pi/512
   m_sin[34]  =  10'b1111010101;     //34pi/512
   m_cos[34]  =  10'b0011111100;     //34pi/512
   m_sin[35]  =  10'b1111010100;     //35pi/512
   m_cos[35]  =  10'b0011111100;     //35pi/512
   m_sin[36]  =  10'b1111010011;     //36pi/512
   m_cos[36]  =  10'b0011111100;     //36pi/512
   m_sin[37]  =  10'b1111010010;     //37pi/512
   m_cos[37]  =  10'b0011111011;     //37pi/512
   m_sin[38]  =  10'b1111010001;     //38pi/512
   m_cos[38]  =  10'b0011111011;     //38pi/512
   m_sin[39]  =  10'b1111001111;     //39pi/512
   m_cos[39]  =  10'b0011111011;     //39pi/512
   m_sin[40]  =  10'b1111001110;     //40pi/512
   m_cos[40]  =  10'b0011111011;     //40pi/512
   m_sin[41]  =  10'b1111001101;     //41pi/512
   m_cos[41]  =  10'b0011111010;     //41pi/512
   m_sin[42]  =  10'b1111001100;     //42pi/512
   m_cos[42]  =  10'b0011111010;     //42pi/512
   m_sin[43]  =  10'b1111001010;     //43pi/512
   m_cos[43]  =  10'b0011111010;     //43pi/512
   m_sin[44]  =  10'b1111001001;     //44pi/512
   m_cos[44]  =  10'b0011111010;     //44pi/512
   m_sin[45]  =  10'b1111001000;     //45pi/512
   m_cos[45]  =  10'b0011111001;     //45pi/512
   m_sin[46]  =  10'b1111000111;     //46pi/512
   m_cos[46]  =  10'b0011111001;     //46pi/512
   m_sin[47]  =  10'b1111000101;     //47pi/512
   m_cos[47]  =  10'b0011111001;     //47pi/512
   m_sin[48]  =  10'b1111000100;     //48pi/512
   m_cos[48]  =  10'b0011111000;     //48pi/512
   m_sin[49]  =  10'b1111000011;     //49pi/512
   m_cos[49]  =  10'b0011111000;     //49pi/512
   m_sin[50]  =  10'b1111000010;     //50pi/512
   m_cos[50]  =  10'b0011111000;     //50pi/512
   m_sin[51]  =  10'b1111000001;     //51pi/512
   m_cos[51]  =  10'b0011111000;     //51pi/512
   m_sin[52]  =  10'b1110111111;     //52pi/512
   m_cos[52]  =  10'b0011110111;     //52pi/512
   m_sin[53]  =  10'b1110111110;     //53pi/512
   m_cos[53]  =  10'b0011110111;     //53pi/512
   m_sin[54]  =  10'b1110111101;     //54pi/512
   m_cos[54]  =  10'b0011110111;     //54pi/512
   m_sin[55]  =  10'b1110111100;     //55pi/512
   m_cos[55]  =  10'b0011110110;     //55pi/512
   m_sin[56]  =  10'b1110111011;     //56pi/512
   m_cos[56]  =  10'b0011110110;     //56pi/512
   m_sin[57]  =  10'b1110111001;     //57pi/512
   m_cos[57]  =  10'b0011110110;     //57pi/512
   m_sin[58]  =  10'b1110111000;     //58pi/512
   m_cos[58]  =  10'b0011110101;     //58pi/512
   m_sin[59]  =  10'b1110110111;     //59pi/512
   m_cos[59]  =  10'b0011110101;     //59pi/512
   m_sin[60]  =  10'b1110110110;     //60pi/512
   m_cos[60]  =  10'b0011110100;     //60pi/512
   m_sin[61]  =  10'b1110110100;     //61pi/512
   m_cos[61]  =  10'b0011110100;     //61pi/512
   m_sin[62]  =  10'b1110110011;     //62pi/512
   m_cos[62]  =  10'b0011110100;     //62pi/512
   m_sin[63]  =  10'b1110110010;     //63pi/512
   m_cos[63]  =  10'b0011110011;     //63pi/512
   m_sin[64]  =  10'b1110110001;     //64pi/512
   m_cos[64]  =  10'b0011110011;     //64pi/512
   m_sin[65]  =  10'b1110110000;     //65pi/512
   m_cos[65]  =  10'b0011110011;     //65pi/512
   m_sin[66]  =  10'b1110101111;     //66pi/512
   m_cos[66]  =  10'b0011110010;     //66pi/512
   m_sin[67]  =  10'b1110101101;     //67pi/512
   m_cos[67]  =  10'b0011110010;     //67pi/512
   m_sin[68]  =  10'b1110101100;     //68pi/512
   m_cos[68]  =  10'b0011110001;     //68pi/512
   m_sin[69]  =  10'b1110101011;     //69pi/512
   m_cos[69]  =  10'b0011110001;     //69pi/512
   m_sin[70]  =  10'b1110101010;     //70pi/512
   m_cos[70]  =  10'b0011110001;     //70pi/512
   m_sin[71]  =  10'b1110101001;     //71pi/512
   m_cos[71]  =  10'b0011110000;     //71pi/512
   m_sin[72]  =  10'b1110100111;     //72pi/512
   m_cos[72]  =  10'b0011110000;     //72pi/512
   m_sin[73]  =  10'b1110100110;     //73pi/512
   m_cos[73]  =  10'b0011101111;     //73pi/512
   m_sin[74]  =  10'b1110100101;     //74pi/512
   m_cos[74]  =  10'b0011101111;     //74pi/512
   m_sin[75]  =  10'b1110100100;     //75pi/512
   m_cos[75]  =  10'b0011101110;     //75pi/512
   m_sin[76]  =  10'b1110100011;     //76pi/512
   m_cos[76]  =  10'b0011101110;     //76pi/512
   m_sin[77]  =  10'b1110100010;     //77pi/512
   m_cos[77]  =  10'b0011101101;     //77pi/512
   m_sin[78]  =  10'b1110100000;     //78pi/512
   m_cos[78]  =  10'b0011101101;     //78pi/512
   m_sin[79]  =  10'b1110011111;     //79pi/512
   m_cos[79]  =  10'b0011101100;     //79pi/512
   m_sin[80]  =  10'b1110011110;     //80pi/512
   m_cos[80]  =  10'b0011101100;     //80pi/512
   m_sin[81]  =  10'b1110011101;     //81pi/512
   m_cos[81]  =  10'b0011101100;     //81pi/512
   m_sin[82]  =  10'b1110011100;     //82pi/512
   m_cos[82]  =  10'b0011101011;     //82pi/512
   m_sin[83]  =  10'b1110011011;     //83pi/512
   m_cos[83]  =  10'b0011101011;     //83pi/512
   m_sin[84]  =  10'b1110011001;     //84pi/512
   m_cos[84]  =  10'b0011101010;     //84pi/512
   m_sin[85]  =  10'b1110011000;     //85pi/512
   m_cos[85]  =  10'b0011101010;     //85pi/512
   m_sin[86]  =  10'b1110010111;     //86pi/512
   m_cos[86]  =  10'b0011101001;     //86pi/512
   m_sin[87]  =  10'b1110010110;     //87pi/512
   m_cos[87]  =  10'b0011101001;     //87pi/512
   m_sin[88]  =  10'b1110010101;     //88pi/512
   m_cos[88]  =  10'b0011101000;     //88pi/512
   m_sin[89]  =  10'b1110010100;     //89pi/512
   m_cos[89]  =  10'b0011100111;     //89pi/512
   m_sin[90]  =  10'b1110010011;     //90pi/512
   m_cos[90]  =  10'b0011100111;     //90pi/512
   m_sin[91]  =  10'b1110010001;     //91pi/512
   m_cos[91]  =  10'b0011100110;     //91pi/512
   m_sin[92]  =  10'b1110010000;     //92pi/512
   m_cos[92]  =  10'b0011100110;     //92pi/512
   m_sin[93]  =  10'b1110001111;     //93pi/512
   m_cos[93]  =  10'b0011100101;     //93pi/512
   m_sin[94]  =  10'b1110001110;     //94pi/512
   m_cos[94]  =  10'b0011100101;     //94pi/512
   m_sin[95]  =  10'b1110001101;     //95pi/512
   m_cos[95]  =  10'b0011100100;     //95pi/512
   m_sin[96]  =  10'b1110001100;     //96pi/512
   m_cos[96]  =  10'b0011100100;     //96pi/512
   m_sin[97]  =  10'b1110001011;     //97pi/512
   m_cos[97]  =  10'b0011100011;     //97pi/512
   m_sin[98]  =  10'b1110001010;     //98pi/512
   m_cos[98]  =  10'b0011100010;     //98pi/512
   m_sin[99]  =  10'b1110001000;     //99pi/512
   m_cos[99]  =  10'b0011100010;     //99pi/512
   m_sin[100]  =  10'b1110000111;     //100pi/512
   m_cos[100]  =  10'b0011100001;     //100pi/512
   m_sin[101]  =  10'b1110000110;     //101pi/512
   m_cos[101]  =  10'b0011100001;     //101pi/512
   m_sin[102]  =  10'b1110000101;     //102pi/512
   m_cos[102]  =  10'b0011100000;     //102pi/512
   m_sin[103]  =  10'b1110000100;     //103pi/512
   m_cos[103]  =  10'b0011011111;     //103pi/512
   m_sin[104]  =  10'b1110000011;     //104pi/512
   m_cos[104]  =  10'b0011011111;     //104pi/512
   m_sin[105]  =  10'b1110000010;     //105pi/512
   m_cos[105]  =  10'b0011011110;     //105pi/512
   m_sin[106]  =  10'b1110000001;     //106pi/512
   m_cos[106]  =  10'b0011011110;     //106pi/512
   m_sin[107]  =  10'b1110000000;     //107pi/512
   m_cos[107]  =  10'b0011011101;     //107pi/512
   m_sin[108]  =  10'b1101111111;     //108pi/512
   m_cos[108]  =  10'b0011011100;     //108pi/512
   m_sin[109]  =  10'b1101111101;     //109pi/512
   m_cos[109]  =  10'b0011011100;     //109pi/512
   m_sin[110]  =  10'b1101111100;     //110pi/512
   m_cos[110]  =  10'b0011011011;     //110pi/512
   m_sin[111]  =  10'b1101111011;     //111pi/512
   m_cos[111]  =  10'b0011011010;     //111pi/512
   m_sin[112]  =  10'b1101111010;     //112pi/512
   m_cos[112]  =  10'b0011011010;     //112pi/512
   m_sin[113]  =  10'b1101111001;     //113pi/512
   m_cos[113]  =  10'b0011011001;     //113pi/512
   m_sin[114]  =  10'b1101111000;     //114pi/512
   m_cos[114]  =  10'b0011011000;     //114pi/512
   m_sin[115]  =  10'b1101110111;     //115pi/512
   m_cos[115]  =  10'b0011011000;     //115pi/512
   m_sin[116]  =  10'b1101110110;     //116pi/512
   m_cos[116]  =  10'b0011010111;     //116pi/512
   m_sin[117]  =  10'b1101110101;     //117pi/512
   m_cos[117]  =  10'b0011010110;     //117pi/512
   m_sin[118]  =  10'b1101110100;     //118pi/512
   m_cos[118]  =  10'b0011010110;     //118pi/512
   m_sin[119]  =  10'b1101110011;     //119pi/512
   m_cos[119]  =  10'b0011010101;     //119pi/512
   m_sin[120]  =  10'b1101110010;     //120pi/512
   m_cos[120]  =  10'b0011010100;     //120pi/512
   m_sin[121]  =  10'b1101110001;     //121pi/512
   m_cos[121]  =  10'b0011010100;     //121pi/512
   m_sin[122]  =  10'b1101110000;     //122pi/512
   m_cos[122]  =  10'b0011010011;     //122pi/512
   m_sin[123]  =  10'b1101101111;     //123pi/512
   m_cos[123]  =  10'b0011010010;     //123pi/512
   m_sin[124]  =  10'b1101101110;     //124pi/512
   m_cos[124]  =  10'b0011010010;     //124pi/512
   m_sin[125]  =  10'b1101101101;     //125pi/512
   m_cos[125]  =  10'b0011010001;     //125pi/512
   m_sin[126]  =  10'b1101101100;     //126pi/512
   m_cos[126]  =  10'b0011010000;     //126pi/512
   m_sin[127]  =  10'b1101101011;     //127pi/512
   m_cos[127]  =  10'b0011001111;     //127pi/512
   m_sin[128]  =  10'b1101101010;     //128pi/512
   m_cos[128]  =  10'b0011001111;     //128pi/512
   m_sin[129]  =  10'b1101101001;     //129pi/512
   m_cos[129]  =  10'b0011001110;     //129pi/512
   m_sin[130]  =  10'b1101101000;     //130pi/512
   m_cos[130]  =  10'b0011001101;     //130pi/512
   m_sin[131]  =  10'b1101100110;     //131pi/512
   m_cos[131]  =  10'b0011001100;     //131pi/512
   m_sin[132]  =  10'b1101100101;     //132pi/512
   m_cos[132]  =  10'b0011001100;     //132pi/512
   m_sin[133]  =  10'b1101100100;     //133pi/512
   m_cos[133]  =  10'b0011001011;     //133pi/512
   m_sin[134]  =  10'b1101100011;     //134pi/512
   m_cos[134]  =  10'b0011001010;     //134pi/512
   m_sin[135]  =  10'b1101100011;     //135pi/512
   m_cos[135]  =  10'b0011001001;     //135pi/512
   m_sin[136]  =  10'b1101100010;     //136pi/512
   m_cos[136]  =  10'b0011001001;     //136pi/512
   m_sin[137]  =  10'b1101100001;     //137pi/512
   m_cos[137]  =  10'b0011001000;     //137pi/512
   m_sin[138]  =  10'b1101100000;     //138pi/512
   m_cos[138]  =  10'b0011000111;     //138pi/512
   m_sin[139]  =  10'b1101011111;     //139pi/512
   m_cos[139]  =  10'b0011000110;     //139pi/512
   m_sin[140]  =  10'b1101011110;     //140pi/512
   m_cos[140]  =  10'b0011000101;     //140pi/512
   m_sin[141]  =  10'b1101011101;     //141pi/512
   m_cos[141]  =  10'b0011000101;     //141pi/512
   m_sin[142]  =  10'b1101011100;     //142pi/512
   m_cos[142]  =  10'b0011000100;     //142pi/512
   m_sin[143]  =  10'b1101011011;     //143pi/512
   m_cos[143]  =  10'b0011000011;     //143pi/512
   m_sin[144]  =  10'b1101011010;     //144pi/512
   m_cos[144]  =  10'b0011000010;     //144pi/512
   m_sin[145]  =  10'b1101011001;     //145pi/512
   m_cos[145]  =  10'b0011000001;     //145pi/512
   m_sin[146]  =  10'b1101011000;     //146pi/512
   m_cos[146]  =  10'b0011000001;     //146pi/512
   m_sin[147]  =  10'b1101010111;     //147pi/512
   m_cos[147]  =  10'b0011000000;     //147pi/512
   m_sin[148]  =  10'b1101010110;     //148pi/512
   m_cos[148]  =  10'b0010111111;     //148pi/512
   m_sin[149]  =  10'b1101010101;     //149pi/512
   m_cos[149]  =  10'b0010111110;     //149pi/512
   m_sin[150]  =  10'b1101010100;     //150pi/512
   m_cos[150]  =  10'b0010111101;     //150pi/512
   m_sin[151]  =  10'b1101010011;     //151pi/512
   m_cos[151]  =  10'b0010111100;     //151pi/512
   m_sin[152]  =  10'b1101010010;     //152pi/512
   m_cos[152]  =  10'b0010111011;     //152pi/512
   m_sin[153]  =  10'b1101010001;     //153pi/512
   m_cos[153]  =  10'b0010111011;     //153pi/512
   m_sin[154]  =  10'b1101010000;     //154pi/512
   m_cos[154]  =  10'b0010111010;     //154pi/512
   m_sin[155]  =  10'b1101001111;     //155pi/512
   m_cos[155]  =  10'b0010111001;     //155pi/512
   m_sin[156]  =  10'b1101001111;     //156pi/512
   m_cos[156]  =  10'b0010111000;     //156pi/512
   m_sin[157]  =  10'b1101001110;     //157pi/512
   m_cos[157]  =  10'b0010110111;     //157pi/512
   m_sin[158]  =  10'b1101001101;     //158pi/512
   m_cos[158]  =  10'b0010110110;     //158pi/512
   m_sin[159]  =  10'b1101001100;     //159pi/512
   m_cos[159]  =  10'b0010110101;     //159pi/512
   m_sin[160]  =  10'b1101001011;     //160pi/512
   m_cos[160]  =  10'b0010110101;     //160pi/512
   m_sin[161]  =  10'b1101001010;     //161pi/512
   m_cos[161]  =  10'b0010110100;     //161pi/512
   m_sin[162]  =  10'b1101001001;     //162pi/512
   m_cos[162]  =  10'b0010110011;     //162pi/512
   m_sin[163]  =  10'b1101001000;     //163pi/512
   m_cos[163]  =  10'b0010110010;     //163pi/512
   m_sin[164]  =  10'b1101000111;     //164pi/512
   m_cos[164]  =  10'b0010110001;     //164pi/512
   m_sin[165]  =  10'b1101000111;     //165pi/512
   m_cos[165]  =  10'b0010110000;     //165pi/512
   m_sin[166]  =  10'b1101000110;     //166pi/512
   m_cos[166]  =  10'b0010101111;     //166pi/512
   m_sin[167]  =  10'b1101000101;     //167pi/512
   m_cos[167]  =  10'b0010101110;     //167pi/512
   m_sin[168]  =  10'b1101000100;     //168pi/512
   m_cos[168]  =  10'b0010101101;     //168pi/512
   m_sin[169]  =  10'b1101000011;     //169pi/512
   m_cos[169]  =  10'b0010101100;     //169pi/512
   m_sin[170]  =  10'b1101000010;     //170pi/512
   m_cos[170]  =  10'b0010101011;     //170pi/512
   m_sin[171]  =  10'b1101000001;     //171pi/512
   m_cos[171]  =  10'b0010101010;     //171pi/512
   m_sin[172]  =  10'b1101000001;     //172pi/512
   m_cos[172]  =  10'b0010101010;     //172pi/512
   m_sin[173]  =  10'b1101000000;     //173pi/512
   m_cos[173]  =  10'b0010101001;     //173pi/512
   m_sin[174]  =  10'b1100111111;     //174pi/512
   m_cos[174]  =  10'b0010101000;     //174pi/512
   m_sin[175]  =  10'b1100111110;     //175pi/512
   m_cos[175]  =  10'b0010100111;     //175pi/512
   m_sin[176]  =  10'b1100111101;     //176pi/512
   m_cos[176]  =  10'b0010100110;     //176pi/512
   m_sin[177]  =  10'b1100111101;     //177pi/512
   m_cos[177]  =  10'b0010100101;     //177pi/512
   m_sin[178]  =  10'b1100111100;     //178pi/512
   m_cos[178]  =  10'b0010100100;     //178pi/512
   m_sin[179]  =  10'b1100111011;     //179pi/512
   m_cos[179]  =  10'b0010100011;     //179pi/512
   m_sin[180]  =  10'b1100111010;     //180pi/512
   m_cos[180]  =  10'b0010100010;     //180pi/512
   m_sin[181]  =  10'b1100111001;     //181pi/512
   m_cos[181]  =  10'b0010100001;     //181pi/512
   m_sin[182]  =  10'b1100111001;     //182pi/512
   m_cos[182]  =  10'b0010100000;     //182pi/512
   m_sin[183]  =  10'b1100111000;     //183pi/512
   m_cos[183]  =  10'b0010011111;     //183pi/512
   m_sin[184]  =  10'b1100110111;     //184pi/512
   m_cos[184]  =  10'b0010011110;     //184pi/512
   m_sin[185]  =  10'b1100110110;     //185pi/512
   m_cos[185]  =  10'b0010011101;     //185pi/512
   m_sin[186]  =  10'b1100110101;     //186pi/512
   m_cos[186]  =  10'b0010011100;     //186pi/512
   m_sin[187]  =  10'b1100110101;     //187pi/512
   m_cos[187]  =  10'b0010011011;     //187pi/512
   m_sin[188]  =  10'b1100110100;     //188pi/512
   m_cos[188]  =  10'b0010011010;     //188pi/512
   m_sin[189]  =  10'b1100110011;     //189pi/512
   m_cos[189]  =  10'b0010011001;     //189pi/512
   m_sin[190]  =  10'b1100110010;     //190pi/512
   m_cos[190]  =  10'b0010011000;     //190pi/512
   m_sin[191]  =  10'b1100110010;     //191pi/512
   m_cos[191]  =  10'b0010010111;     //191pi/512
   m_sin[192]  =  10'b1100110001;     //192pi/512
   m_cos[192]  =  10'b0010010110;     //192pi/512
   m_sin[193]  =  10'b1100110000;     //193pi/512
   m_cos[193]  =  10'b0010010101;     //193pi/512
   m_sin[194]  =  10'b1100101111;     //194pi/512
   m_cos[194]  =  10'b0010010100;     //194pi/512
   m_sin[195]  =  10'b1100101111;     //195pi/512
   m_cos[195]  =  10'b0010010011;     //195pi/512
   m_sin[196]  =  10'b1100101110;     //196pi/512
   m_cos[196]  =  10'b0010010010;     //196pi/512
   m_sin[197]  =  10'b1100101101;     //197pi/512
   m_cos[197]  =  10'b0010010001;     //197pi/512
   m_sin[198]  =  10'b1100101101;     //198pi/512
   m_cos[198]  =  10'b0010010000;     //198pi/512
   m_sin[199]  =  10'b1100101100;     //199pi/512
   m_cos[199]  =  10'b0010001111;     //199pi/512
   m_sin[200]  =  10'b1100101011;     //200pi/512
   m_cos[200]  =  10'b0010001110;     //200pi/512
   m_sin[201]  =  10'b1100101010;     //201pi/512
   m_cos[201]  =  10'b0010001101;     //201pi/512
   m_sin[202]  =  10'b1100101010;     //202pi/512
   m_cos[202]  =  10'b0010001100;     //202pi/512
   m_sin[203]  =  10'b1100101001;     //203pi/512
   m_cos[203]  =  10'b0010001011;     //203pi/512
   m_sin[204]  =  10'b1100101000;     //204pi/512
   m_cos[204]  =  10'b0010001010;     //204pi/512
   m_sin[205]  =  10'b1100101000;     //205pi/512
   m_cos[205]  =  10'b0010001000;     //205pi/512
   m_sin[206]  =  10'b1100100111;     //206pi/512
   m_cos[206]  =  10'b0010000111;     //206pi/512
   m_sin[207]  =  10'b1100100110;     //207pi/512
   m_cos[207]  =  10'b0010000110;     //207pi/512
   m_sin[208]  =  10'b1100100110;     //208pi/512
   m_cos[208]  =  10'b0010000101;     //208pi/512
   m_sin[209]  =  10'b1100100101;     //209pi/512
   m_cos[209]  =  10'b0010000100;     //209pi/512
   m_sin[210]  =  10'b1100100100;     //210pi/512
   m_cos[210]  =  10'b0010000011;     //210pi/512
   m_sin[211]  =  10'b1100100100;     //211pi/512
   m_cos[211]  =  10'b0010000010;     //211pi/512
   m_sin[212]  =  10'b1100100011;     //212pi/512
   m_cos[212]  =  10'b0010000001;     //212pi/512
   m_sin[213]  =  10'b1100100011;     //213pi/512
   m_cos[213]  =  10'b0010000000;     //213pi/512
   m_sin[214]  =  10'b1100100010;     //214pi/512
   m_cos[214]  =  10'b0001111111;     //214pi/512
   m_sin[215]  =  10'b1100100001;     //215pi/512
   m_cos[215]  =  10'b0001111110;     //215pi/512
   m_sin[216]  =  10'b1100100001;     //216pi/512
   m_cos[216]  =  10'b0001111101;     //216pi/512
   m_sin[217]  =  10'b1100100000;     //217pi/512
   m_cos[217]  =  10'b0001111011;     //217pi/512
   m_sin[218]  =  10'b1100011111;     //218pi/512
   m_cos[218]  =  10'b0001111010;     //218pi/512
   m_sin[219]  =  10'b1100011111;     //219pi/512
   m_cos[219]  =  10'b0001111001;     //219pi/512
   m_sin[220]  =  10'b1100011110;     //220pi/512
   m_cos[220]  =  10'b0001111000;     //220pi/512
   m_sin[221]  =  10'b1100011110;     //221pi/512
   m_cos[221]  =  10'b0001110111;     //221pi/512
   m_sin[222]  =  10'b1100011101;     //222pi/512
   m_cos[222]  =  10'b0001110110;     //222pi/512
   m_sin[223]  =  10'b1100011100;     //223pi/512
   m_cos[223]  =  10'b0001110101;     //223pi/512
   m_sin[224]  =  10'b1100011100;     //224pi/512
   m_cos[224]  =  10'b0001110100;     //224pi/512
   m_sin[225]  =  10'b1100011011;     //225pi/512
   m_cos[225]  =  10'b0001110011;     //225pi/512
   m_sin[226]  =  10'b1100011011;     //226pi/512
   m_cos[226]  =  10'b0001110001;     //226pi/512
   m_sin[227]  =  10'b1100011010;     //227pi/512
   m_cos[227]  =  10'b0001110000;     //227pi/512
   m_sin[228]  =  10'b1100011010;     //228pi/512
   m_cos[228]  =  10'b0001101111;     //228pi/512
   m_sin[229]  =  10'b1100011001;     //229pi/512
   m_cos[229]  =  10'b0001101110;     //229pi/512
   m_sin[230]  =  10'b1100011001;     //230pi/512
   m_cos[230]  =  10'b0001101101;     //230pi/512
   m_sin[231]  =  10'b1100011000;     //231pi/512
   m_cos[231]  =  10'b0001101100;     //231pi/512
   m_sin[232]  =  10'b1100011000;     //232pi/512
   m_cos[232]  =  10'b0001101011;     //232pi/512
   m_sin[233]  =  10'b1100010111;     //233pi/512
   m_cos[233]  =  10'b0001101010;     //233pi/512
   m_sin[234]  =  10'b1100010110;     //234pi/512
   m_cos[234]  =  10'b0001101000;     //234pi/512
   m_sin[235]  =  10'b1100010110;     //235pi/512
   m_cos[235]  =  10'b0001100111;     //235pi/512
   m_sin[236]  =  10'b1100010101;     //236pi/512
   m_cos[236]  =  10'b0001100110;     //236pi/512
   m_sin[237]  =  10'b1100010101;     //237pi/512
   m_cos[237]  =  10'b0001100101;     //237pi/512
   m_sin[238]  =  10'b1100010100;     //238pi/512
   m_cos[238]  =  10'b0001100100;     //238pi/512
   m_sin[239]  =  10'b1100010100;     //239pi/512
   m_cos[239]  =  10'b0001100011;     //239pi/512
   m_sin[240]  =  10'b1100010011;     //240pi/512
   m_cos[240]  =  10'b0001100001;     //240pi/512
   m_sin[241]  =  10'b1100010011;     //241pi/512
   m_cos[241]  =  10'b0001100000;     //241pi/512
   m_sin[242]  =  10'b1100010011;     //242pi/512
   m_cos[242]  =  10'b0001011111;     //242pi/512
   m_sin[243]  =  10'b1100010010;     //243pi/512
   m_cos[243]  =  10'b0001011110;     //243pi/512
   m_sin[244]  =  10'b1100010010;     //244pi/512
   m_cos[244]  =  10'b0001011101;     //244pi/512
   m_sin[245]  =  10'b1100010001;     //245pi/512
   m_cos[245]  =  10'b0001011100;     //245pi/512
   m_sin[246]  =  10'b1100010001;     //246pi/512
   m_cos[246]  =  10'b0001011010;     //246pi/512
   m_sin[247]  =  10'b1100010000;     //247pi/512
   m_cos[247]  =  10'b0001011001;     //247pi/512
   m_sin[248]  =  10'b1100010000;     //248pi/512
   m_cos[248]  =  10'b0001011000;     //248pi/512
   m_sin[249]  =  10'b1100001111;     //249pi/512
   m_cos[249]  =  10'b0001010111;     //249pi/512
   m_sin[250]  =  10'b1100001111;     //250pi/512
   m_cos[250]  =  10'b0001010110;     //250pi/512
   m_sin[251]  =  10'b1100001111;     //251pi/512
   m_cos[251]  =  10'b0001010101;     //251pi/512
   m_sin[252]  =  10'b1100001110;     //252pi/512
   m_cos[252]  =  10'b0001010011;     //252pi/512
   m_sin[253]  =  10'b1100001110;     //253pi/512
   m_cos[253]  =  10'b0001010010;     //253pi/512
   m_sin[254]  =  10'b1100001101;     //254pi/512
   m_cos[254]  =  10'b0001010001;     //254pi/512
   m_sin[255]  =  10'b1100001101;     //255pi/512
   m_cos[255]  =  10'b0001010000;     //255pi/512
   m_sin[256]  =  10'b1100001101;     //256pi/512
   m_cos[256]  =  10'b0001001111;     //256pi/512
   m_sin[257]  =  10'b1100001100;     //257pi/512
   m_cos[257]  =  10'b0001001101;     //257pi/512
   m_sin[258]  =  10'b1100001100;     //258pi/512
   m_cos[258]  =  10'b0001001100;     //258pi/512
   m_sin[259]  =  10'b1100001011;     //259pi/512
   m_cos[259]  =  10'b0001001011;     //259pi/512
   m_sin[260]  =  10'b1100001011;     //260pi/512
   m_cos[260]  =  10'b0001001010;     //260pi/512
   m_sin[261]  =  10'b1100001011;     //261pi/512
   m_cos[261]  =  10'b0001001001;     //261pi/512
   m_sin[262]  =  10'b1100001010;     //262pi/512
   m_cos[262]  =  10'b0001000111;     //262pi/512
   m_sin[263]  =  10'b1100001010;     //263pi/512
   m_cos[263]  =  10'b0001000110;     //263pi/512
   m_sin[264]  =  10'b1100001010;     //264pi/512
   m_cos[264]  =  10'b0001000101;     //264pi/512
   m_sin[265]  =  10'b1100001001;     //265pi/512
   m_cos[265]  =  10'b0001000100;     //265pi/512
   m_sin[266]  =  10'b1100001001;     //266pi/512
   m_cos[266]  =  10'b0001000011;     //266pi/512
   m_sin[267]  =  10'b1100001001;     //267pi/512
   m_cos[267]  =  10'b0001000001;     //267pi/512
   m_sin[268]  =  10'b1100001000;     //268pi/512
   m_cos[268]  =  10'b0001000000;     //268pi/512
   m_sin[269]  =  10'b1100001000;     //269pi/512
   m_cos[269]  =  10'b0000111111;     //269pi/512
   m_sin[270]  =  10'b1100001000;     //270pi/512
   m_cos[270]  =  10'b0000111110;     //270pi/512
   m_sin[271]  =  10'b1100000111;     //271pi/512
   m_cos[271]  =  10'b0000111100;     //271pi/512
   m_sin[272]  =  10'b1100000111;     //272pi/512
   m_cos[272]  =  10'b0000111011;     //272pi/512
   m_sin[273]  =  10'b1100000111;     //273pi/512
   m_cos[273]  =  10'b0000111010;     //273pi/512
   m_sin[274]  =  10'b1100000110;     //274pi/512
   m_cos[274]  =  10'b0000111001;     //274pi/512
   m_sin[275]  =  10'b1100000110;     //275pi/512
   m_cos[275]  =  10'b0000111000;     //275pi/512
   m_sin[276]  =  10'b1100000110;     //276pi/512
   m_cos[276]  =  10'b0000110110;     //276pi/512
   m_sin[277]  =  10'b1100000110;     //277pi/512
   m_cos[277]  =  10'b0000110101;     //277pi/512
   m_sin[278]  =  10'b1100000101;     //278pi/512
   m_cos[278]  =  10'b0000110100;     //278pi/512
   m_sin[279]  =  10'b1100000101;     //279pi/512
   m_cos[279]  =  10'b0000110011;     //279pi/512
   m_sin[280]  =  10'b1100000101;     //280pi/512
   m_cos[280]  =  10'b0000110001;     //280pi/512
   m_sin[281]  =  10'b1100000101;     //281pi/512
   m_cos[281]  =  10'b0000110000;     //281pi/512
   m_sin[282]  =  10'b1100000100;     //282pi/512
   m_cos[282]  =  10'b0000101111;     //282pi/512
   m_sin[283]  =  10'b1100000100;     //283pi/512
   m_cos[283]  =  10'b0000101110;     //283pi/512
   m_sin[284]  =  10'b1100000100;     //284pi/512
   m_cos[284]  =  10'b0000101101;     //284pi/512
   m_sin[285]  =  10'b1100000100;     //285pi/512
   m_cos[285]  =  10'b0000101011;     //285pi/512
   m_sin[286]  =  10'b1100000100;     //286pi/512
   m_cos[286]  =  10'b0000101010;     //286pi/512
   m_sin[287]  =  10'b1100000011;     //287pi/512
   m_cos[287]  =  10'b0000101001;     //287pi/512
   m_sin[288]  =  10'b1100000011;     //288pi/512
   m_cos[288]  =  10'b0000101000;     //288pi/512
   m_sin[289]  =  10'b1100000011;     //289pi/512
   m_cos[289]  =  10'b0000100110;     //289pi/512
   m_sin[290]  =  10'b1100000011;     //290pi/512
   m_cos[290]  =  10'b0000100101;     //290pi/512
   m_sin[291]  =  10'b1100000011;     //291pi/512
   m_cos[291]  =  10'b0000100100;     //291pi/512
   m_sin[292]  =  10'b1100000010;     //292pi/512
   m_cos[292]  =  10'b0000100011;     //292pi/512
   m_sin[293]  =  10'b1100000010;     //293pi/512
   m_cos[293]  =  10'b0000100001;     //293pi/512
   m_sin[294]  =  10'b1100000010;     //294pi/512
   m_cos[294]  =  10'b0000100000;     //294pi/512
   m_sin[295]  =  10'b1100000010;     //295pi/512
   m_cos[295]  =  10'b0000011111;     //295pi/512
   m_sin[296]  =  10'b1100000010;     //296pi/512
   m_cos[296]  =  10'b0000011110;     //296pi/512
   m_sin[297]  =  10'b1100000010;     //297pi/512
   m_cos[297]  =  10'b0000011100;     //297pi/512
   m_sin[298]  =  10'b1100000001;     //298pi/512
   m_cos[298]  =  10'b0000011011;     //298pi/512
   m_sin[299]  =  10'b1100000001;     //299pi/512
   m_cos[299]  =  10'b0000011010;     //299pi/512
   m_sin[300]  =  10'b1100000001;     //300pi/512
   m_cos[300]  =  10'b0000011001;     //300pi/512
   m_sin[301]  =  10'b1100000001;     //301pi/512
   m_cos[301]  =  10'b0000010111;     //301pi/512
   m_sin[302]  =  10'b1100000001;     //302pi/512
   m_cos[302]  =  10'b0000010110;     //302pi/512
   m_sin[303]  =  10'b1100000001;     //303pi/512
   m_cos[303]  =  10'b0000010101;     //303pi/512
   m_sin[304]  =  10'b1100000001;     //304pi/512
   m_cos[304]  =  10'b0000010100;     //304pi/512
   m_sin[305]  =  10'b1100000001;     //305pi/512
   m_cos[305]  =  10'b0000010010;     //305pi/512
   m_sin[306]  =  10'b1100000001;     //306pi/512
   m_cos[306]  =  10'b0000010001;     //306pi/512
   m_sin[307]  =  10'b1100000001;     //307pi/512
   m_cos[307]  =  10'b0000010000;     //307pi/512
   m_sin[308]  =  10'b1100000000;     //308pi/512
   m_cos[308]  =  10'b0000001111;     //308pi/512
   m_sin[309]  =  10'b1100000000;     //309pi/512
   m_cos[309]  =  10'b0000001101;     //309pi/512
   m_sin[310]  =  10'b1100000000;     //310pi/512
   m_cos[310]  =  10'b0000001100;     //310pi/512
   m_sin[311]  =  10'b1100000000;     //311pi/512
   m_cos[311]  =  10'b0000001011;     //311pi/512
   m_sin[312]  =  10'b1100000000;     //312pi/512
   m_cos[312]  =  10'b0000001010;     //312pi/512
   m_sin[313]  =  10'b1100000000;     //313pi/512
   m_cos[313]  =  10'b0000001000;     //313pi/512
   m_sin[314]  =  10'b1100000000;     //314pi/512
   m_cos[314]  =  10'b0000000111;     //314pi/512
   m_sin[315]  =  10'b1100000000;     //315pi/512
   m_cos[315]  =  10'b0000000110;     //315pi/512
   m_sin[316]  =  10'b1100000000;     //316pi/512
   m_cos[316]  =  10'b0000000101;     //316pi/512
   m_sin[317]  =  10'b1100000000;     //317pi/512
   m_cos[317]  =  10'b0000000011;     //317pi/512
   m_sin[318]  =  10'b1100000000;     //318pi/512
   m_cos[318]  =  10'b0000000010;     //318pi/512
   m_sin[319]  =  10'b1100000000;     //319pi/512
   m_cos[319]  =  10'b0000000001;     //319pi/512
   m_sin[320]  =  10'b1100000000;     //320pi/512
   m_cos[320]  =  10'b0000000000;     //320pi/512
   m_sin[321]  =  10'b1100000000;     //321pi/512
   m_cos[321]  =  10'b1111111111;     //321pi/512
   m_sin[322]  =  10'b1100000000;     //322pi/512
   m_cos[322]  =  10'b1111111101;     //322pi/512
   m_sin[323]  =  10'b1100000000;     //323pi/512
   m_cos[323]  =  10'b1111111100;     //323pi/512
   m_sin[324]  =  10'b1100000000;     //324pi/512
   m_cos[324]  =  10'b1111111011;     //324pi/512
   m_sin[325]  =  10'b1100000000;     //325pi/512
   m_cos[325]  =  10'b1111111010;     //325pi/512
   m_sin[326]  =  10'b1100000000;     //326pi/512
   m_cos[326]  =  10'b1111111000;     //326pi/512
   m_sin[327]  =  10'b1100000000;     //327pi/512
   m_cos[327]  =  10'b1111110111;     //327pi/512
   m_sin[328]  =  10'b1100000000;     //328pi/512
   m_cos[328]  =  10'b1111110110;     //328pi/512
   m_sin[329]  =  10'b1100000000;     //329pi/512
   m_cos[329]  =  10'b1111110101;     //329pi/512
   m_sin[330]  =  10'b1100000000;     //330pi/512
   m_cos[330]  =  10'b1111110011;     //330pi/512
   m_sin[331]  =  10'b1100000000;     //331pi/512
   m_cos[331]  =  10'b1111110010;     //331pi/512
   m_sin[332]  =  10'b1100000000;     //332pi/512
   m_cos[332]  =  10'b1111110001;     //332pi/512
   m_sin[333]  =  10'b1100000001;     //333pi/512
   m_cos[333]  =  10'b1111110000;     //333pi/512
   m_sin[334]  =  10'b1100000001;     //334pi/512
   m_cos[334]  =  10'b1111101110;     //334pi/512
   m_sin[335]  =  10'b1100000001;     //335pi/512
   m_cos[335]  =  10'b1111101101;     //335pi/512
   m_sin[336]  =  10'b1100000001;     //336pi/512
   m_cos[336]  =  10'b1111101100;     //336pi/512
   m_sin[337]  =  10'b1100000001;     //337pi/512
   m_cos[337]  =  10'b1111101011;     //337pi/512
   m_sin[338]  =  10'b1100000001;     //338pi/512
   m_cos[338]  =  10'b1111101001;     //338pi/512
   m_sin[339]  =  10'b1100000001;     //339pi/512
   m_cos[339]  =  10'b1111101000;     //339pi/512
   m_sin[340]  =  10'b1100000001;     //340pi/512
   m_cos[340]  =  10'b1111100111;     //340pi/512
   m_sin[341]  =  10'b1100000001;     //341pi/512
   m_cos[341]  =  10'b1111100110;     //341pi/512
   m_sin[342]  =  10'b1100000001;     //342pi/512
   m_cos[342]  =  10'b1111100100;     //342pi/512
   m_sin[343]  =  10'b1100000010;     //343pi/512
   m_cos[343]  =  10'b1111100011;     //343pi/512
   m_sin[344]  =  10'b1100000010;     //344pi/512
   m_cos[344]  =  10'b1111100010;     //344pi/512
   m_sin[345]  =  10'b1100000010;     //345pi/512
   m_cos[345]  =  10'b1111100001;     //345pi/512
   m_sin[346]  =  10'b1100000010;     //346pi/512
   m_cos[346]  =  10'b1111011111;     //346pi/512
   m_sin[347]  =  10'b1100000010;     //347pi/512
   m_cos[347]  =  10'b1111011110;     //347pi/512
   m_sin[348]  =  10'b1100000010;     //348pi/512
   m_cos[348]  =  10'b1111011101;     //348pi/512
   m_sin[349]  =  10'b1100000011;     //349pi/512
   m_cos[349]  =  10'b1111011100;     //349pi/512
   m_sin[350]  =  10'b1100000011;     //350pi/512
   m_cos[350]  =  10'b1111011010;     //350pi/512
   m_sin[351]  =  10'b1100000011;     //351pi/512
   m_cos[351]  =  10'b1111011001;     //351pi/512
   m_sin[352]  =  10'b1100000011;     //352pi/512
   m_cos[352]  =  10'b1111011000;     //352pi/512
   m_sin[353]  =  10'b1100000011;     //353pi/512
   m_cos[353]  =  10'b1111010111;     //353pi/512
   m_sin[354]  =  10'b1100000100;     //354pi/512
   m_cos[354]  =  10'b1111010101;     //354pi/512
   m_sin[355]  =  10'b1100000100;     //355pi/512
   m_cos[355]  =  10'b1111010100;     //355pi/512
   m_sin[356]  =  10'b1100000100;     //356pi/512
   m_cos[356]  =  10'b1111010011;     //356pi/512
   m_sin[357]  =  10'b1100000100;     //357pi/512
   m_cos[357]  =  10'b1111010010;     //357pi/512
   m_sin[358]  =  10'b1100000100;     //358pi/512
   m_cos[358]  =  10'b1111010001;     //358pi/512
   m_sin[359]  =  10'b1100000101;     //359pi/512
   m_cos[359]  =  10'b1111001111;     //359pi/512
   m_sin[360]  =  10'b1100000101;     //360pi/512
   m_cos[360]  =  10'b1111001110;     //360pi/512
   m_sin[361]  =  10'b1100000101;     //361pi/512
   m_cos[361]  =  10'b1111001101;     //361pi/512
   m_sin[362]  =  10'b1100000101;     //362pi/512
   m_cos[362]  =  10'b1111001100;     //362pi/512
   m_sin[363]  =  10'b1100000110;     //363pi/512
   m_cos[363]  =  10'b1111001010;     //363pi/512
   m_sin[364]  =  10'b1100000110;     //364pi/512
   m_cos[364]  =  10'b1111001001;     //364pi/512
   m_sin[365]  =  10'b1100000110;     //365pi/512
   m_cos[365]  =  10'b1111001000;     //365pi/512
   m_sin[366]  =  10'b1100000110;     //366pi/512
   m_cos[366]  =  10'b1111000111;     //366pi/512
   m_sin[367]  =  10'b1100000111;     //367pi/512
   m_cos[367]  =  10'b1111000101;     //367pi/512
   m_sin[368]  =  10'b1100000111;     //368pi/512
   m_cos[368]  =  10'b1111000100;     //368pi/512
   m_sin[369]  =  10'b1100000111;     //369pi/512
   m_cos[369]  =  10'b1111000011;     //369pi/512
   m_sin[370]  =  10'b1100001000;     //370pi/512
   m_cos[370]  =  10'b1111000010;     //370pi/512
   m_sin[371]  =  10'b1100001000;     //371pi/512
   m_cos[371]  =  10'b1111000001;     //371pi/512
   m_sin[372]  =  10'b1100001000;     //372pi/512
   m_cos[372]  =  10'b1110111111;     //372pi/512
   m_sin[373]  =  10'b1100001001;     //373pi/512
   m_cos[373]  =  10'b1110111110;     //373pi/512
   m_sin[374]  =  10'b1100001001;     //374pi/512
   m_cos[374]  =  10'b1110111101;     //374pi/512
   m_sin[375]  =  10'b1100001001;     //375pi/512
   m_cos[375]  =  10'b1110111100;     //375pi/512
   m_sin[376]  =  10'b1100001010;     //376pi/512
   m_cos[376]  =  10'b1110111011;     //376pi/512
   m_sin[377]  =  10'b1100001010;     //377pi/512
   m_cos[377]  =  10'b1110111001;     //377pi/512
   m_sin[378]  =  10'b1100001010;     //378pi/512
   m_cos[378]  =  10'b1110111000;     //378pi/512
   m_sin[379]  =  10'b1100001011;     //379pi/512
   m_cos[379]  =  10'b1110110111;     //379pi/512
   m_sin[380]  =  10'b1100001011;     //380pi/512
   m_cos[380]  =  10'b1110110110;     //380pi/512
   m_sin[381]  =  10'b1100001011;     //381pi/512
   m_cos[381]  =  10'b1110110100;     //381pi/512
   m_sin[382]  =  10'b1100001100;     //382pi/512
   m_cos[382]  =  10'b1110110011;     //382pi/512
   m_sin[383]  =  10'b1100001100;     //383pi/512
   m_cos[383]  =  10'b1110110010;     //383pi/512
   m_sin[384]  =  10'b1100001101;     //384pi/512
   m_cos[384]  =  10'b1110110001;     //384pi/512
   m_sin[385]  =  10'b1100001101;     //385pi/512
   m_cos[385]  =  10'b1110110000;     //385pi/512
   m_sin[386]  =  10'b1100001101;     //386pi/512
   m_cos[386]  =  10'b1110101111;     //386pi/512
   m_sin[387]  =  10'b1100001110;     //387pi/512
   m_cos[387]  =  10'b1110101101;     //387pi/512
   m_sin[388]  =  10'b1100001110;     //388pi/512
   m_cos[388]  =  10'b1110101100;     //388pi/512
   m_sin[389]  =  10'b1100001111;     //389pi/512
   m_cos[389]  =  10'b1110101011;     //389pi/512
   m_sin[390]  =  10'b1100001111;     //390pi/512
   m_cos[390]  =  10'b1110101010;     //390pi/512
   m_sin[391]  =  10'b1100001111;     //391pi/512
   m_cos[391]  =  10'b1110101001;     //391pi/512
   m_sin[392]  =  10'b1100010000;     //392pi/512
   m_cos[392]  =  10'b1110100111;     //392pi/512
   m_sin[393]  =  10'b1100010000;     //393pi/512
   m_cos[393]  =  10'b1110100110;     //393pi/512
   m_sin[394]  =  10'b1100010001;     //394pi/512
   m_cos[394]  =  10'b1110100101;     //394pi/512
   m_sin[395]  =  10'b1100010001;     //395pi/512
   m_cos[395]  =  10'b1110100100;     //395pi/512
   m_sin[396]  =  10'b1100010010;     //396pi/512
   m_cos[396]  =  10'b1110100011;     //396pi/512
   m_sin[397]  =  10'b1100010010;     //397pi/512
   m_cos[397]  =  10'b1110100010;     //397pi/512
   m_sin[398]  =  10'b1100010011;     //398pi/512
   m_cos[398]  =  10'b1110100000;     //398pi/512
   m_sin[399]  =  10'b1100010011;     //399pi/512
   m_cos[399]  =  10'b1110011111;     //399pi/512
   m_sin[400]  =  10'b1100010011;     //400pi/512
   m_cos[400]  =  10'b1110011110;     //400pi/512
   m_sin[401]  =  10'b1100010100;     //401pi/512
   m_cos[401]  =  10'b1110011101;     //401pi/512
   m_sin[402]  =  10'b1100010100;     //402pi/512
   m_cos[402]  =  10'b1110011100;     //402pi/512
   m_sin[403]  =  10'b1100010101;     //403pi/512
   m_cos[403]  =  10'b1110011011;     //403pi/512
   m_sin[404]  =  10'b1100010101;     //404pi/512
   m_cos[404]  =  10'b1110011001;     //404pi/512
   m_sin[405]  =  10'b1100010110;     //405pi/512
   m_cos[405]  =  10'b1110011000;     //405pi/512
   m_sin[406]  =  10'b1100010110;     //406pi/512
   m_cos[406]  =  10'b1110010111;     //406pi/512
   m_sin[407]  =  10'b1100010111;     //407pi/512
   m_cos[407]  =  10'b1110010110;     //407pi/512
   m_sin[408]  =  10'b1100011000;     //408pi/512
   m_cos[408]  =  10'b1110010101;     //408pi/512
   m_sin[409]  =  10'b1100011000;     //409pi/512
   m_cos[409]  =  10'b1110010100;     //409pi/512
   m_sin[410]  =  10'b1100011001;     //410pi/512
   m_cos[410]  =  10'b1110010011;     //410pi/512
   m_sin[411]  =  10'b1100011001;     //411pi/512
   m_cos[411]  =  10'b1110010001;     //411pi/512
   m_sin[412]  =  10'b1100011010;     //412pi/512
   m_cos[412]  =  10'b1110010000;     //412pi/512
   m_sin[413]  =  10'b1100011010;     //413pi/512
   m_cos[413]  =  10'b1110001111;     //413pi/512
   m_sin[414]  =  10'b1100011011;     //414pi/512
   m_cos[414]  =  10'b1110001110;     //414pi/512
   m_sin[415]  =  10'b1100011011;     //415pi/512
   m_cos[415]  =  10'b1110001101;     //415pi/512
   m_sin[416]  =  10'b1100011100;     //416pi/512
   m_cos[416]  =  10'b1110001100;     //416pi/512
   m_sin[417]  =  10'b1100011100;     //417pi/512
   m_cos[417]  =  10'b1110001011;     //417pi/512
   m_sin[418]  =  10'b1100011101;     //418pi/512
   m_cos[418]  =  10'b1110001010;     //418pi/512
   m_sin[419]  =  10'b1100011110;     //419pi/512
   m_cos[419]  =  10'b1110001000;     //419pi/512
   m_sin[420]  =  10'b1100011110;     //420pi/512
   m_cos[420]  =  10'b1110000111;     //420pi/512
   m_sin[421]  =  10'b1100011111;     //421pi/512
   m_cos[421]  =  10'b1110000110;     //421pi/512
   m_sin[422]  =  10'b1100011111;     //422pi/512
   m_cos[422]  =  10'b1110000101;     //422pi/512
   m_sin[423]  =  10'b1100100000;     //423pi/512
   m_cos[423]  =  10'b1110000100;     //423pi/512
   m_sin[424]  =  10'b1100100001;     //424pi/512
   m_cos[424]  =  10'b1110000011;     //424pi/512
   m_sin[425]  =  10'b1100100001;     //425pi/512
   m_cos[425]  =  10'b1110000010;     //425pi/512
   m_sin[426]  =  10'b1100100010;     //426pi/512
   m_cos[426]  =  10'b1110000001;     //426pi/512
   m_sin[427]  =  10'b1100100011;     //427pi/512
   m_cos[427]  =  10'b1110000000;     //427pi/512
   m_sin[428]  =  10'b1100100011;     //428pi/512
   m_cos[428]  =  10'b1101111111;     //428pi/512
   m_sin[429]  =  10'b1100100100;     //429pi/512
   m_cos[429]  =  10'b1101111101;     //429pi/512
   m_sin[430]  =  10'b1100100100;     //430pi/512
   m_cos[430]  =  10'b1101111100;     //430pi/512
   m_sin[431]  =  10'b1100100101;     //431pi/512
   m_cos[431]  =  10'b1101111011;     //431pi/512
   m_sin[432]  =  10'b1100100110;     //432pi/512
   m_cos[432]  =  10'b1101111010;     //432pi/512
   m_sin[433]  =  10'b1100100110;     //433pi/512
   m_cos[433]  =  10'b1101111001;     //433pi/512
   m_sin[434]  =  10'b1100100111;     //434pi/512
   m_cos[434]  =  10'b1101111000;     //434pi/512
   m_sin[435]  =  10'b1100101000;     //435pi/512
   m_cos[435]  =  10'b1101110111;     //435pi/512
   m_sin[436]  =  10'b1100101000;     //436pi/512
   m_cos[436]  =  10'b1101110110;     //436pi/512
   m_sin[437]  =  10'b1100101001;     //437pi/512
   m_cos[437]  =  10'b1101110101;     //437pi/512
   m_sin[438]  =  10'b1100101010;     //438pi/512
   m_cos[438]  =  10'b1101110100;     //438pi/512
   m_sin[439]  =  10'b1100101010;     //439pi/512
   m_cos[439]  =  10'b1101110011;     //439pi/512
   m_sin[440]  =  10'b1100101011;     //440pi/512
   m_cos[440]  =  10'b1101110010;     //440pi/512
   m_sin[441]  =  10'b1100101100;     //441pi/512
   m_cos[441]  =  10'b1101110001;     //441pi/512
   m_sin[442]  =  10'b1100101101;     //442pi/512
   m_cos[442]  =  10'b1101110000;     //442pi/512
   m_sin[443]  =  10'b1100101101;     //443pi/512
   m_cos[443]  =  10'b1101101111;     //443pi/512
   m_sin[444]  =  10'b1100101110;     //444pi/512
   m_cos[444]  =  10'b1101101110;     //444pi/512
   m_sin[445]  =  10'b1100101111;     //445pi/512
   m_cos[445]  =  10'b1101101101;     //445pi/512
   m_sin[446]  =  10'b1100101111;     //446pi/512
   m_cos[446]  =  10'b1101101100;     //446pi/512
   m_sin[447]  =  10'b1100110000;     //447pi/512
   m_cos[447]  =  10'b1101101011;     //447pi/512
   m_sin[448]  =  10'b1100110001;     //448pi/512
   m_cos[448]  =  10'b1101101010;     //448pi/512
   m_sin[449]  =  10'b1100110010;     //449pi/512
   m_cos[449]  =  10'b1101101001;     //449pi/512
   m_sin[450]  =  10'b1100110010;     //450pi/512
   m_cos[450]  =  10'b1101101000;     //450pi/512
   m_sin[451]  =  10'b1100110011;     //451pi/512
   m_cos[451]  =  10'b1101100110;     //451pi/512
   m_sin[452]  =  10'b1100110100;     //452pi/512
   m_cos[452]  =  10'b1101100101;     //452pi/512
   m_sin[453]  =  10'b1100110101;     //453pi/512
   m_cos[453]  =  10'b1101100100;     //453pi/512
   m_sin[454]  =  10'b1100110101;     //454pi/512
   m_cos[454]  =  10'b1101100011;     //454pi/512
   m_sin[455]  =  10'b1100110110;     //455pi/512
   m_cos[455]  =  10'b1101100011;     //455pi/512
   m_sin[456]  =  10'b1100110111;     //456pi/512
   m_cos[456]  =  10'b1101100010;     //456pi/512
   m_sin[457]  =  10'b1100111000;     //457pi/512
   m_cos[457]  =  10'b1101100001;     //457pi/512
   m_sin[458]  =  10'b1100111001;     //458pi/512
   m_cos[458]  =  10'b1101100000;     //458pi/512
   m_sin[459]  =  10'b1100111001;     //459pi/512
   m_cos[459]  =  10'b1101011111;     //459pi/512
   m_sin[460]  =  10'b1100111010;     //460pi/512
   m_cos[460]  =  10'b1101011110;     //460pi/512
   m_sin[461]  =  10'b1100111011;     //461pi/512
   m_cos[461]  =  10'b1101011101;     //461pi/512
   m_sin[462]  =  10'b1100111100;     //462pi/512
   m_cos[462]  =  10'b1101011100;     //462pi/512
   m_sin[463]  =  10'b1100111101;     //463pi/512
   m_cos[463]  =  10'b1101011011;     //463pi/512
   m_sin[464]  =  10'b1100111101;     //464pi/512
   m_cos[464]  =  10'b1101011010;     //464pi/512
   m_sin[465]  =  10'b1100111110;     //465pi/512
   m_cos[465]  =  10'b1101011001;     //465pi/512
   m_sin[466]  =  10'b1100111111;     //466pi/512
   m_cos[466]  =  10'b1101011000;     //466pi/512
   m_sin[467]  =  10'b1101000000;     //467pi/512
   m_cos[467]  =  10'b1101010111;     //467pi/512
   m_sin[468]  =  10'b1101000001;     //468pi/512
   m_cos[468]  =  10'b1101010110;     //468pi/512
   m_sin[469]  =  10'b1101000001;     //469pi/512
   m_cos[469]  =  10'b1101010101;     //469pi/512
   m_sin[470]  =  10'b1101000010;     //470pi/512
   m_cos[470]  =  10'b1101010100;     //470pi/512
   m_sin[471]  =  10'b1101000011;     //471pi/512
   m_cos[471]  =  10'b1101010011;     //471pi/512
   m_sin[472]  =  10'b1101000100;     //472pi/512
   m_cos[472]  =  10'b1101010010;     //472pi/512
   m_sin[473]  =  10'b1101000101;     //473pi/512
   m_cos[473]  =  10'b1101010001;     //473pi/512
   m_sin[474]  =  10'b1101000110;     //474pi/512
   m_cos[474]  =  10'b1101010000;     //474pi/512
   m_sin[475]  =  10'b1101000111;     //475pi/512
   m_cos[475]  =  10'b1101001111;     //475pi/512
   m_sin[476]  =  10'b1101000111;     //476pi/512
   m_cos[476]  =  10'b1101001111;     //476pi/512
   m_sin[477]  =  10'b1101001000;     //477pi/512
   m_cos[477]  =  10'b1101001110;     //477pi/512
   m_sin[478]  =  10'b1101001001;     //478pi/512
   m_cos[478]  =  10'b1101001101;     //478pi/512
   m_sin[479]  =  10'b1101001010;     //479pi/512
   m_cos[479]  =  10'b1101001100;     //479pi/512
   m_sin[480]  =  10'b1101001011;     //480pi/512
   m_cos[480]  =  10'b1101001011;     //480pi/512
   m_sin[481]  =  10'b1101001100;     //481pi/512
   m_cos[481]  =  10'b1101001010;     //481pi/512
   m_sin[482]  =  10'b1101001101;     //482pi/512
   m_cos[482]  =  10'b1101001001;     //482pi/512
   m_sin[483]  =  10'b1101001110;     //483pi/512
   m_cos[483]  =  10'b1101001000;     //483pi/512
   m_sin[484]  =  10'b1101001111;     //484pi/512
   m_cos[484]  =  10'b1101000111;     //484pi/512
   m_sin[485]  =  10'b1101001111;     //485pi/512
   m_cos[485]  =  10'b1101000111;     //485pi/512
   m_sin[486]  =  10'b1101010000;     //486pi/512
   m_cos[486]  =  10'b1101000110;     //486pi/512
   m_sin[487]  =  10'b1101010001;     //487pi/512
   m_cos[487]  =  10'b1101000101;     //487pi/512
   m_sin[488]  =  10'b1101010010;     //488pi/512
   m_cos[488]  =  10'b1101000100;     //488pi/512
   m_sin[489]  =  10'b1101010011;     //489pi/512
   m_cos[489]  =  10'b1101000011;     //489pi/512
   m_sin[490]  =  10'b1101010100;     //490pi/512
   m_cos[490]  =  10'b1101000010;     //490pi/512
   m_sin[491]  =  10'b1101010101;     //491pi/512
   m_cos[491]  =  10'b1101000001;     //491pi/512
   m_sin[492]  =  10'b1101010110;     //492pi/512
   m_cos[492]  =  10'b1101000001;     //492pi/512
   m_sin[493]  =  10'b1101010111;     //493pi/512
   m_cos[493]  =  10'b1101000000;     //493pi/512
   m_sin[494]  =  10'b1101011000;     //494pi/512
   m_cos[494]  =  10'b1100111111;     //494pi/512
   m_sin[495]  =  10'b1101011001;     //495pi/512
   m_cos[495]  =  10'b1100111110;     //495pi/512
   m_sin[496]  =  10'b1101011010;     //496pi/512
   m_cos[496]  =  10'b1100111101;     //496pi/512
   m_sin[497]  =  10'b1101011011;     //497pi/512
   m_cos[497]  =  10'b1100111101;     //497pi/512
   m_sin[498]  =  10'b1101011100;     //498pi/512
   m_cos[498]  =  10'b1100111100;     //498pi/512
   m_sin[499]  =  10'b1101011101;     //499pi/512
   m_cos[499]  =  10'b1100111011;     //499pi/512
   m_sin[500]  =  10'b1101011110;     //500pi/512
   m_cos[500]  =  10'b1100111010;     //500pi/512
   m_sin[501]  =  10'b1101011111;     //501pi/512
   m_cos[501]  =  10'b1100111001;     //501pi/512
   m_sin[502]  =  10'b1101100000;     //502pi/512
   m_cos[502]  =  10'b1100111001;     //502pi/512
   m_sin[503]  =  10'b1101100001;     //503pi/512
   m_cos[503]  =  10'b1100111000;     //503pi/512
   m_sin[504]  =  10'b1101100010;     //504pi/512
   m_cos[504]  =  10'b1100110111;     //504pi/512
   m_sin[505]  =  10'b1101100011;     //505pi/512
   m_cos[505]  =  10'b1100110110;     //505pi/512
   m_sin[506]  =  10'b1101100011;     //506pi/512
   m_cos[506]  =  10'b1100110101;     //506pi/512
   m_sin[507]  =  10'b1101100100;     //507pi/512
   m_cos[507]  =  10'b1100110101;     //507pi/512
   m_sin[508]  =  10'b1101100101;     //508pi/512
   m_cos[508]  =  10'b1100110100;     //508pi/512
   m_sin[509]  =  10'b1101100110;     //509pi/512
   m_cos[509]  =  10'b1100110011;     //509pi/512
   m_sin[510]  =  10'b1101101000;     //510pi/512
   m_cos[510]  =  10'b1100110010;     //510pi/512
   m_sin[511]  =  10'b1101101001;     //511pi/512
   m_cos[511]  =  10'b1100110010;     //511pi/512
end
endmodule