module  TWIDLE_14_bit_STAGE1  #(parameter N = 256, SIZE = 8, bit_width_tw = 14) (
    input                               clk,
    input          [SIZE        -2:0]   rd_ptr_angle,
    input                               en, 

    output reg signed [bit_width_tw-1:0]   cos_data,
    output reg signed [bit_width_tw-1:0]   sin_data
 );

reg signed [bit_width_tw-1:0]  cos  [127:0];
reg signed [bit_width_tw-1:0]  sin  [127:0];

localparam  coefficient =  $clog2(256/N);

wire [6:0] rd_ptr = rd_ptr_angle << coefficient;

always @(posedge clk) begin
  if (en) begin
    cos_data <= cos [rd_ptr];
    sin_data <= sin [rd_ptr];
  end
end


initial begin

   sin[0]  =  14'b00000000000000;     //0pi/256
   cos[0]  =  14'b01000000000000;     //0pi/256
   sin[1]  =  14'b11111110011011;     //2pi/256
   cos[1]  =  14'b00111111111110;     //2pi/256
   sin[2]  =  14'b11111100110111;     //4pi/256
   cos[2]  =  14'b00111111111011;     //4pi/256
   sin[3]  =  14'b11111011010011;     //6pi/256
   cos[3]  =  14'b00111111110100;     //6pi/256
   sin[4]  =  14'b11111001101111;     //8pi/256
   cos[4]  =  14'b00111111101100;     //8pi/256
   sin[5]  =  14'b11111000001011;     //10pi/256
   cos[5]  =  14'b00111111100001;     //10pi/256
   sin[6]  =  14'b11110110100111;     //12pi/256
   cos[6]  =  14'b00111111010011;     //12pi/256
   sin[7]  =  14'b11110101000100;     //14pi/256
   cos[7]  =  14'b00111111000011;     //14pi/256
   sin[8]  =  14'b11110011100001;     //16pi/256
   cos[8]  =  14'b00111110110001;     //16pi/256
   sin[9]  =  14'b11110001111111;     //18pi/256
   cos[9]  =  14'b00111110011100;     //18pi/256
   sin[10]  =  14'b11110000011101;     //20pi/256
   cos[10]  =  14'b00111110000101;     //20pi/256
   sin[11]  =  14'b11101110111100;     //22pi/256
   cos[11]  =  14'b00111101101011;     //22pi/256
   sin[12]  =  14'b11101101011011;     //24pi/256
   cos[12]  =  14'b00111101001111;     //24pi/256
   sin[13]  =  14'b11101011111011;     //26pi/256
   cos[13]  =  14'b00111100110001;     //26pi/256
   sin[14]  =  14'b11101010011100;     //28pi/256
   cos[14]  =  14'b00111100010000;     //28pi/256
   sin[15]  =  14'b11101000111110;     //30pi/256
   cos[15]  =  14'b00111011101101;     //30pi/256
   sin[16]  =  14'b11100111100001;     //32pi/256
   cos[16]  =  14'b00111011001000;     //32pi/256
   sin[17]  =  14'b11100110000100;     //34pi/256
   cos[17]  =  14'b00111010100000;     //34pi/256
   sin[18]  =  14'b11100100101001;     //36pi/256
   cos[18]  =  14'b00111001110110;     //36pi/256
   sin[19]  =  14'b11100011001110;     //38pi/256
   cos[19]  =  14'b00111001001010;     //38pi/256
   sin[20]  =  14'b11100001110101;     //40pi/256
   cos[20]  =  14'b00111000011100;     //40pi/256
   sin[21]  =  14'b11100000011101;     //42pi/256
   cos[21]  =  14'b00110111101011;     //42pi/256
   sin[22]  =  14'b11011111000110;     //44pi/256
   cos[22]  =  14'b00110110111001;     //44pi/256
   sin[23]  =  14'b11011101110001;     //46pi/256
   cos[23]  =  14'b00110110000100;     //46pi/256
   sin[24]  =  14'b11011100011100;     //48pi/256
   cos[24]  =  14'b00110101001101;     //48pi/256
   sin[25]  =  14'b11011011001001;     //50pi/256
   cos[25]  =  14'b00110100010100;     //50pi/256
   sin[26]  =  14'b11011001111000;     //52pi/256
   cos[26]  =  14'b00110011011001;     //52pi/256
   sin[27]  =  14'b11011000101000;     //54pi/256
   cos[27]  =  14'b00110010011101;     //54pi/256
   sin[28]  =  14'b11010111011010;     //56pi/256
   cos[28]  =  14'b00110001011110;     //56pi/256
   sin[29]  =  14'b11010110001101;     //58pi/256
   cos[29]  =  14'b00110000011101;     //58pi/256
   sin[30]  =  14'b11010101000001;     //60pi/256
   cos[30]  =  14'b00101111011010;     //60pi/256
   sin[31]  =  14'b11010011111000;     //62pi/256
   cos[31]  =  14'b00101110010110;     //62pi/256
   sin[32]  =  14'b11010010110000;     //64pi/256
   cos[32]  =  14'b00101101010000;     //64pi/256
   sin[33]  =  14'b11010001101001;     //66pi/256
   cos[33]  =  14'b00101100001000;     //66pi/256
   sin[34]  =  14'b11010000100101;     //68pi/256
   cos[34]  =  14'b00101010111110;     //68pi/256
   sin[35]  =  14'b11001111100010;     //70pi/256
   cos[35]  =  14'b00101001110011;     //70pi/256
   sin[36]  =  14'b11001110100010;     //72pi/256
   cos[36]  =  14'b00101000100110;     //72pi/256
   sin[37]  =  14'b11001101100011;     //74pi/256
   cos[37]  =  14'b00100111010111;     //74pi/256
   sin[38]  =  14'b11001100100110;     //76pi/256
   cos[38]  =  14'b00100110000111;     //76pi/256
   sin[39]  =  14'b11001011101011;     //78pi/256
   cos[39]  =  14'b00100100110110;     //78pi/256
   sin[40]  =  14'b11001010110010;     //80pi/256
   cos[40]  =  14'b00100011100011;     //80pi/256
   sin[41]  =  14'b11001001111011;     //82pi/256
   cos[41]  =  14'b00100010001111;     //82pi/256
   sin[42]  =  14'b11001001000111;     //84pi/256
   cos[42]  =  14'b00100000111001;     //84pi/256
   sin[43]  =  14'b11001000010100;     //86pi/256
   cos[43]  =  14'b00011111100010;     //86pi/256
   sin[44]  =  14'b11000111100100;     //88pi/256
   cos[44]  =  14'b00011110001010;     //88pi/256
   sin[45]  =  14'b11000110110101;     //90pi/256
   cos[45]  =  14'b00011100110001;     //90pi/256
   sin[46]  =  14'b11000110001001;     //92pi/256
   cos[46]  =  14'b00011011010111;     //92pi/256
   sin[47]  =  14'b11000101011111;     //94pi/256
   cos[47]  =  14'b00011001111011;     //94pi/256
   sin[48]  =  14'b11000100111000;     //96pi/256
   cos[48]  =  14'b00011000011111;     //96pi/256
   sin[49]  =  14'b11000100010010;     //98pi/256
   cos[49]  =  14'b00010111000010;     //98pi/256
   sin[50]  =  14'b11000011101111;     //100pi/256
   cos[50]  =  14'b00010101100011;     //100pi/256
   sin[51]  =  14'b11000011001111;     //102pi/256
   cos[51]  =  14'b00010100000100;     //102pi/256
   sin[52]  =  14'b11000010110000;     //104pi/256
   cos[52]  =  14'b00010010100101;     //104pi/256
   sin[53]  =  14'b11000010010100;     //106pi/256
   cos[53]  =  14'b00010001000100;     //106pi/256
   sin[54]  =  14'b11000001111011;     //108pi/256
   cos[54]  =  14'b00001111100011;     //108pi/256
   sin[55]  =  14'b11000001100100;     //110pi/256
   cos[55]  =  14'b00001110000001;     //110pi/256
   sin[56]  =  14'b11000001001111;     //112pi/256
   cos[56]  =  14'b00001100011111;     //112pi/256
   sin[57]  =  14'b11000000111100;     //114pi/256
   cos[57]  =  14'b00001010111100;     //114pi/256
   sin[58]  =  14'b11000000101100;     //116pi/256
   cos[58]  =  14'b00001001011001;     //116pi/256
   sin[59]  =  14'b11000000011111;     //118pi/256
   cos[59]  =  14'b00000111110101;     //118pi/256
   sin[60]  =  14'b11000000010100;     //120pi/256
   cos[60]  =  14'b00000110010001;     //120pi/256
   sin[61]  =  14'b11000000001011;     //122pi/256
   cos[61]  =  14'b00000100101101;     //122pi/256
   sin[62]  =  14'b11000000000101;     //124pi/256
   cos[62]  =  14'b00000011001000;     //124pi/256
   sin[63]  =  14'b11000000000001;     //126pi/256
   cos[63]  =  14'b00000001100100;     //126pi/256
   sin[64]  =  14'b11000000000000;     //128pi/256
   cos[64]  =  14'b00000000000000;     //128pi/256
   sin[65]  =  14'b11000000000001;     //130pi/256
   cos[65]  =  14'b11111110011011;     //130pi/256
   sin[66]  =  14'b11000000000101;     //132pi/256
   cos[66]  =  14'b11111100110111;     //132pi/256
   sin[67]  =  14'b11000000001011;     //134pi/256
   cos[67]  =  14'b11111011010011;     //134pi/256
   sin[68]  =  14'b11000000010100;     //136pi/256
   cos[68]  =  14'b11111001101111;     //136pi/256
   sin[69]  =  14'b11000000011111;     //138pi/256
   cos[69]  =  14'b11111000001011;     //138pi/256
   sin[70]  =  14'b11000000101100;     //140pi/256
   cos[70]  =  14'b11110110100111;     //140pi/256
   sin[71]  =  14'b11000000111100;     //142pi/256
   cos[71]  =  14'b11110101000100;     //142pi/256
   sin[72]  =  14'b11000001001111;     //144pi/256
   cos[72]  =  14'b11110011100001;     //144pi/256
   sin[73]  =  14'b11000001100100;     //146pi/256
   cos[73]  =  14'b11110001111111;     //146pi/256
   sin[74]  =  14'b11000001111011;     //148pi/256
   cos[74]  =  14'b11110000011101;     //148pi/256
   sin[75]  =  14'b11000010010100;     //150pi/256
   cos[75]  =  14'b11101110111100;     //150pi/256
   sin[76]  =  14'b11000010110000;     //152pi/256
   cos[76]  =  14'b11101101011011;     //152pi/256
   sin[77]  =  14'b11000011001111;     //154pi/256
   cos[77]  =  14'b11101011111011;     //154pi/256
   sin[78]  =  14'b11000011101111;     //156pi/256
   cos[78]  =  14'b11101010011100;     //156pi/256
   sin[79]  =  14'b11000100010010;     //158pi/256
   cos[79]  =  14'b11101000111110;     //158pi/256
   sin[80]  =  14'b11000100111000;     //160pi/256
   cos[80]  =  14'b11100111100001;     //160pi/256
   sin[81]  =  14'b11000101011111;     //162pi/256
   cos[81]  =  14'b11100110000100;     //162pi/256
   sin[82]  =  14'b11000110001001;     //164pi/256
   cos[82]  =  14'b11100100101001;     //164pi/256
   sin[83]  =  14'b11000110110101;     //166pi/256
   cos[83]  =  14'b11100011001110;     //166pi/256
   sin[84]  =  14'b11000111100100;     //168pi/256
   cos[84]  =  14'b11100001110101;     //168pi/256
   sin[85]  =  14'b11001000010100;     //170pi/256
   cos[85]  =  14'b11100000011101;     //170pi/256
   sin[86]  =  14'b11001001000111;     //172pi/256
   cos[86]  =  14'b11011111000110;     //172pi/256
   sin[87]  =  14'b11001001111011;     //174pi/256
   cos[87]  =  14'b11011101110001;     //174pi/256
   sin[88]  =  14'b11001010110010;     //176pi/256
   cos[88]  =  14'b11011100011100;     //176pi/256
   sin[89]  =  14'b11001011101011;     //178pi/256
   cos[89]  =  14'b11011011001001;     //178pi/256
   sin[90]  =  14'b11001100100110;     //180pi/256
   cos[90]  =  14'b11011001111000;     //180pi/256
   sin[91]  =  14'b11001101100011;     //182pi/256
   cos[91]  =  14'b11011000101000;     //182pi/256
   sin[92]  =  14'b11001110100010;     //184pi/256
   cos[92]  =  14'b11010111011010;     //184pi/256
   sin[93]  =  14'b11001111100010;     //186pi/256
   cos[93]  =  14'b11010110001101;     //186pi/256
   sin[94]  =  14'b11010000100101;     //188pi/256
   cos[94]  =  14'b11010101000001;     //188pi/256
   sin[95]  =  14'b11010001101001;     //190pi/256
   cos[95]  =  14'b11010011111000;     //190pi/256
   sin[96]  =  14'b11010010110000;     //192pi/256
   cos[96]  =  14'b11010010110000;     //192pi/256
   sin[97]  =  14'b11010011111000;     //194pi/256
   cos[97]  =  14'b11010001101001;     //194pi/256
   sin[98]  =  14'b11010101000001;     //196pi/256
   cos[98]  =  14'b11010000100101;     //196pi/256
   sin[99]  =  14'b11010110001101;     //198pi/256
   cos[99]  =  14'b11001111100010;     //198pi/256
   sin[100]  =  14'b11010111011010;     //200pi/256
   cos[100]  =  14'b11001110100010;     //200pi/256
   sin[101]  =  14'b11011000101000;     //202pi/256
   cos[101]  =  14'b11001101100011;     //202pi/256
   sin[102]  =  14'b11011001111000;     //204pi/256
   cos[102]  =  14'b11001100100110;     //204pi/256
   sin[103]  =  14'b11011011001001;     //206pi/256
   cos[103]  =  14'b11001011101011;     //206pi/256
   sin[104]  =  14'b11011100011100;     //208pi/256
   cos[104]  =  14'b11001010110010;     //208pi/256
   sin[105]  =  14'b11011101110001;     //210pi/256
   cos[105]  =  14'b11001001111011;     //210pi/256
   sin[106]  =  14'b11011111000110;     //212pi/256
   cos[106]  =  14'b11001001000111;     //212pi/256
   sin[107]  =  14'b11100000011101;     //214pi/256
   cos[107]  =  14'b11001000010100;     //214pi/256
   sin[108]  =  14'b11100001110101;     //216pi/256
   cos[108]  =  14'b11000111100100;     //216pi/256
   sin[109]  =  14'b11100011001110;     //218pi/256
   cos[109]  =  14'b11000110110101;     //218pi/256
   sin[110]  =  14'b11100100101001;     //220pi/256
   cos[110]  =  14'b11000110001001;     //220pi/256
   sin[111]  =  14'b11100110000100;     //222pi/256
   cos[111]  =  14'b11000101011111;     //222pi/256
   sin[112]  =  14'b11100111100001;     //224pi/256
   cos[112]  =  14'b11000100111000;     //224pi/256
   sin[113]  =  14'b11101000111110;     //226pi/256
   cos[113]  =  14'b11000100010010;     //226pi/256
   sin[114]  =  14'b11101010011100;     //228pi/256
   cos[114]  =  14'b11000011101111;     //228pi/256
   sin[115]  =  14'b11101011111011;     //230pi/256
   cos[115]  =  14'b11000011001111;     //230pi/256
   sin[116]  =  14'b11101101011011;     //232pi/256
   cos[116]  =  14'b11000010110000;     //232pi/256
   sin[117]  =  14'b11101110111100;     //234pi/256
   cos[117]  =  14'b11000010010100;     //234pi/256
   sin[118]  =  14'b11110000011101;     //236pi/256
   cos[118]  =  14'b11000001111011;     //236pi/256
   sin[119]  =  14'b11110001111111;     //238pi/256
   cos[119]  =  14'b11000001100100;     //238pi/256
   sin[120]  =  14'b11110011100001;     //240pi/256
   cos[120]  =  14'b11000001001111;     //240pi/256
   sin[121]  =  14'b11110101000100;     //242pi/256
   cos[121]  =  14'b11000000111100;     //242pi/256
   sin[122]  =  14'b11110110100111;     //244pi/256
   cos[122]  =  14'b11000000101100;     //244pi/256
   sin[123]  =  14'b11111000001011;     //246pi/256
   cos[123]  =  14'b11000000011111;     //246pi/256
   sin[124]  =  14'b11111001101111;     //248pi/256
   cos[124]  =  14'b11000000010100;     //248pi/256
   sin[125]  =  14'b11111011010011;     //250pi/256
   cos[125]  =  14'b11000000001011;     //250pi/256
   sin[126]  =  14'b11111100110111;     //252pi/256
   cos[126]  =  14'b11000000000101;     //252pi/256
   sin[127]  =  14'b11111110011011;     //254pi/256
   cos[127]  =  14'b11000000000001;     //254pi/256

end
endmodule