
module  TWIDLE_14_bit_STAGE2  #(parameter N = 256, SIZE = 8, bit_width_tw = 14) (
    input                               clk,
    input          [SIZE        -3:0]   rd_ptr_angle,
    input                               en, 

    output  reg signed [bit_width_tw-1:0]   cos_data,
    output  reg signed [bit_width_tw-1:0]   sin_data
 );

reg signed [bit_width_tw-1:0]  cos  [64:0];
reg signed [bit_width_tw-1:0]  sin  [64:0];

localparam  coefficient =  $clog2(256/N);

wire [6:0] rd_ptr = rd_ptr_angle << coefficient;

always @(posedge clk) begin
  if (en) begin
    cos_data <= cos [rd_ptr];
    sin_data <= sin [rd_ptr];
  end
end


initial begin
   sin[0]  =  14'b00000000000000;     //0pi/256
   cos[0]  =  14'b01000000000000;     //0pi/256
   sin[1]  =  14'b11111100110111;     //4pi/256
   cos[1]  =  14'b00111111111011;     //4pi/256
   sin[2]  =  14'b11111001101111;     //8pi/256
   cos[2]  =  14'b00111111101100;     //8pi/256
   sin[3]  =  14'b11110110100111;     //12pi/256
   cos[3]  =  14'b00111111010011;     //12pi/256
   sin[4]  =  14'b11110011100001;     //16pi/256
   cos[4]  =  14'b00111110110001;     //16pi/256
   sin[5]  =  14'b11110000011101;     //20pi/256
   cos[5]  =  14'b00111110000101;     //20pi/256
   sin[6]  =  14'b11101101011011;     //24pi/256
   cos[6]  =  14'b00111101001111;     //24pi/256
   sin[7]  =  14'b11101010011100;     //28pi/256
   cos[7]  =  14'b00111100010000;     //28pi/256
   sin[8]  =  14'b11100111100001;     //32pi/256
   cos[8]  =  14'b00111011001000;     //32pi/256
   sin[9]  =  14'b11100100101001;     //36pi/256
   cos[9]  =  14'b00111001110110;     //36pi/256
   sin[10]  =  14'b11100001110101;     //40pi/256
   cos[10]  =  14'b00111000011100;     //40pi/256
   sin[11]  =  14'b11011111000110;     //44pi/256
   cos[11]  =  14'b00110110111001;     //44pi/256
   sin[12]  =  14'b11011100011100;     //48pi/256
   cos[12]  =  14'b00110101001101;     //48pi/256
   sin[13]  =  14'b11011001111000;     //52pi/256
   cos[13]  =  14'b00110011011001;     //52pi/256
   sin[14]  =  14'b11010111011010;     //56pi/256
   cos[14]  =  14'b00110001011110;     //56pi/256
   sin[15]  =  14'b11010101000001;     //60pi/256
   cos[15]  =  14'b00101111011010;     //60pi/256
   sin[16]  =  14'b11010010110000;     //64pi/256
   cos[16]  =  14'b00101101010000;     //64pi/256
   sin[17]  =  14'b11010000100101;     //68pi/256
   cos[17]  =  14'b00101010111110;     //68pi/256
   sin[18]  =  14'b11001110100010;     //72pi/256
   cos[18]  =  14'b00101000100110;     //72pi/256
   sin[19]  =  14'b11001100100110;     //76pi/256
   cos[19]  =  14'b00100110000111;     //76pi/256
   sin[20]  =  14'b11001010110010;     //80pi/256
   cos[20]  =  14'b00100011100011;     //80pi/256
   sin[21]  =  14'b11001001000111;     //84pi/256
   cos[21]  =  14'b00100000111001;     //84pi/256
   sin[22]  =  14'b11000111100100;     //88pi/256
   cos[22]  =  14'b00011110001010;     //88pi/256
   sin[23]  =  14'b11000110001001;     //92pi/256
   cos[23]  =  14'b00011011010111;     //92pi/256
   sin[24]  =  14'b11000100111000;     //96pi/256
   cos[24]  =  14'b00011000011111;     //96pi/256
   sin[25]  =  14'b11000011101111;     //100pi/256
   cos[25]  =  14'b00010101100011;     //100pi/256
   sin[26]  =  14'b11000010110000;     //104pi/256
   cos[26]  =  14'b00010010100101;     //104pi/256
   sin[27]  =  14'b11000001111011;     //108pi/256
   cos[27]  =  14'b00001111100011;     //108pi/256
   sin[28]  =  14'b11000001001111;     //112pi/256
   cos[28]  =  14'b00001100011111;     //112pi/256
   sin[29]  =  14'b11000000101100;     //116pi/256
   cos[29]  =  14'b00001001011001;     //116pi/256
   sin[30]  =  14'b11000000010100;     //120pi/256
   cos[30]  =  14'b00000110010001;     //120pi/256
   sin[31]  =  14'b11000000000101;     //124pi/256
   cos[31]  =  14'b00000011001000;     //124pi/256
   sin[32]  =  14'b11000000000000;     //128pi/256
   cos[32]  =  14'b00000000000000;     //128pi/256
   sin[33]  =  14'b11000000000101;     //132pi/256
   cos[33]  =  14'b11111100110111;     //132pi/256
   sin[34]  =  14'b11000000010100;     //136pi/256
   cos[34]  =  14'b11111001101111;     //136pi/256
   sin[35]  =  14'b11000000101100;     //140pi/256
   cos[35]  =  14'b11110110100111;     //140pi/256
   sin[36]  =  14'b11000001001111;     //144pi/256
   cos[36]  =  14'b11110011100001;     //144pi/256
   sin[37]  =  14'b11000001111011;     //148pi/256
   cos[37]  =  14'b11110000011101;     //148pi/256
   sin[38]  =  14'b11000010110000;     //152pi/256
   cos[38]  =  14'b11101101011011;     //152pi/256
   sin[39]  =  14'b11000011101111;     //156pi/256
   cos[39]  =  14'b11101010011100;     //156pi/256
   sin[40]  =  14'b11000100111000;     //160pi/256
   cos[40]  =  14'b11100111100001;     //160pi/256
   sin[41]  =  14'b11000110001001;     //164pi/256
   cos[41]  =  14'b11100100101001;     //164pi/256
   sin[42]  =  14'b11000111100100;     //168pi/256
   cos[42]  =  14'b11100001110101;     //168pi/256
   sin[43]  =  14'b11001001000111;     //172pi/256
   cos[43]  =  14'b11011111000110;     //172pi/256
   sin[44]  =  14'b11001010110010;     //176pi/256
   cos[44]  =  14'b11011100011100;     //176pi/256
   sin[45]  =  14'b11001100100110;     //180pi/256
   cos[45]  =  14'b11011001111000;     //180pi/256
   sin[46]  =  14'b11001110100010;     //184pi/256
   cos[46]  =  14'b11010111011010;     //184pi/256
   sin[47]  =  14'b11010000100101;     //188pi/256
   cos[47]  =  14'b11010101000001;     //188pi/256
   sin[48]  =  14'b11010010110000;     //192pi/256
   cos[48]  =  14'b11010010110000;     //192pi/256
   sin[49]  =  14'b11010101000001;     //196pi/256
   cos[49]  =  14'b11010000100101;     //196pi/256
   sin[50]  =  14'b11010111011010;     //200pi/256
   cos[50]  =  14'b11001110100010;     //200pi/256
   sin[51]  =  14'b11011001111000;     //204pi/256
   cos[51]  =  14'b11001100100110;     //204pi/256
   sin[52]  =  14'b11011100011100;     //208pi/256
   cos[52]  =  14'b11001010110010;     //208pi/256
   sin[53]  =  14'b11011111000110;     //212pi/256
   cos[53]  =  14'b11001001000111;     //212pi/256
   sin[54]  =  14'b11100001110101;     //216pi/256
   cos[54]  =  14'b11000111100100;     //216pi/256
   sin[55]  =  14'b11100100101001;     //220pi/256
   cos[55]  =  14'b11000110001001;     //220pi/256
   sin[56]  =  14'b11100111100001;     //224pi/256
   cos[56]  =  14'b11000100111000;     //224pi/256
   sin[57]  =  14'b11101010011100;     //228pi/256
   cos[57]  =  14'b11000011101111;     //228pi/256
   sin[58]  =  14'b11101101011011;     //232pi/256
   cos[58]  =  14'b11000010110000;     //232pi/256
   sin[59]  =  14'b11110000011101;     //236pi/256
   cos[59]  =  14'b11000001111011;     //236pi/256
   sin[60]  =  14'b11110011100001;     //240pi/256
   cos[60]  =  14'b11000001001111;     //240pi/256
   sin[61]  =  14'b11110110100111;     //244pi/256
   cos[61]  =  14'b11000000101100;     //244pi/256
   sin[62]  =  14'b11111001101111;     //248pi/256
   cos[62]  =  14'b11000000010100;     //248pi/256
   sin[63]  =  14'b11111100110111;     //252pi/256
   cos[63]  =  14'b11000000000101;     //252pi/256
end

endmodule