module  M_TWIDLE_16_B_0_5_v  #(parameter SIZE = 10, word_length_tw = 16) (
    input            clk,
    input            en_rd,
    input   [10:0]   rd_ptr_angle,
    input            en_modf,
    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );
reg signed [word_length_tw-1:0]  cos    [511:0];
reg signed [word_length_tw-1:0]  sin    [511:0];
reg signed [word_length_tw-1:0]  m_cos  [511:0];
reg signed [word_length_tw-1:0]  m_sin  [511:0];
reg signed [word_length_tw-1:0]  cos_temp;
reg signed [word_length_tw-1:0]  sin_temp;
reg signed [word_length_tw-1:0]  m_cos_temp;
reg signed [word_length_tw-1:0]  m_sin_temp;
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & ~ en_modf) begin
                  cos_temp           <= cos   [rd_ptr_angle];
                  sin_temp           <= sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & en_modf) begin
                  m_cos_temp           <= m_cos   [rd_ptr_angle];
                  m_sin_temp           <= m_sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(*) begin 
             if (en_modf) begin
                  cos_data           <= m_cos_temp;
                  sin_data           <= m_sin_temp;
             end else begin
                  cos_data           <= cos_temp;
                  sin_data           <= sin_temp;
             end 
        end
initial begin
   sin[0]  =  16'b0000000000000000;     //0pi/512
   cos[0]  =  16'b0100000000000000;     //0pi/512
   sin[1]  =  16'b1111111110011011;     //1pi/512
   cos[1]  =  16'b0011111111111111;     //1pi/512
   sin[2]  =  16'b1111111100110111;     //2pi/512
   cos[2]  =  16'b0011111111111110;     //2pi/512
   sin[3]  =  16'b1111111011010010;     //3pi/512
   cos[3]  =  16'b0011111111111101;     //3pi/512
   sin[4]  =  16'b1111111001101110;     //4pi/512
   cos[4]  =  16'b0011111111111011;     //4pi/512
   sin[5]  =  16'b1111111000001001;     //5pi/512
   cos[5]  =  16'b0011111111111000;     //5pi/512
   sin[6]  =  16'b1111110110100101;     //6pi/512
   cos[6]  =  16'b0011111111110100;     //6pi/512
   sin[7]  =  16'b1111110101000000;     //7pi/512
   cos[7]  =  16'b0011111111110000;     //7pi/512
   sin[8]  =  16'b1111110011011100;     //8pi/512
   cos[8]  =  16'b0011111111101100;     //8pi/512
   sin[9]  =  16'b1111110001111000;     //9pi/512
   cos[9]  =  16'b0011111111100111;     //9pi/512
   sin[10]  =  16'b1111110000010011;     //10pi/512
   cos[10]  =  16'b0011111111100001;     //10pi/512
   sin[11]  =  16'b1111101110101111;     //11pi/512
   cos[11]  =  16'b0011111111011010;     //11pi/512
   sin[12]  =  16'b1111101101001011;     //12pi/512
   cos[12]  =  16'b0011111111010011;     //12pi/512
   sin[13]  =  16'b1111101011100110;     //13pi/512
   cos[13]  =  16'b0011111111001011;     //13pi/512
   sin[14]  =  16'b1111101010000010;     //14pi/512
   cos[14]  =  16'b0011111111000011;     //14pi/512
   sin[15]  =  16'b1111101000011110;     //15pi/512
   cos[15]  =  16'b0011111110111010;     //15pi/512
   sin[16]  =  16'b1111100110111010;     //16pi/512
   cos[16]  =  16'b0011111110110001;     //16pi/512
   sin[17]  =  16'b1111100101010110;     //17pi/512
   cos[17]  =  16'b0011111110100110;     //17pi/512
   sin[18]  =  16'b1111100011110010;     //18pi/512
   cos[18]  =  16'b0011111110011100;     //18pi/512
   sin[19]  =  16'b1111100010001110;     //19pi/512
   cos[19]  =  16'b0011111110010000;     //19pi/512
   sin[20]  =  16'b1111100000101010;     //20pi/512
   cos[20]  =  16'b0011111110000100;     //20pi/512
   sin[21]  =  16'b1111011111000111;     //21pi/512
   cos[21]  =  16'b0011111101111000;     //21pi/512
   sin[22]  =  16'b1111011101100011;     //22pi/512
   cos[22]  =  16'b0011111101101010;     //22pi/512
   sin[23]  =  16'b1111011011111111;     //23pi/512
   cos[23]  =  16'b0011111101011101;     //23pi/512
   sin[24]  =  16'b1111011010011100;     //24pi/512
   cos[24]  =  16'b0011111101001110;     //24pi/512
   sin[25]  =  16'b1111011000111001;     //25pi/512
   cos[25]  =  16'b0011111100111111;     //25pi/512
   sin[26]  =  16'b1111010111010101;     //26pi/512
   cos[26]  =  16'b0011111100101111;     //26pi/512
   sin[27]  =  16'b1111010101110010;     //27pi/512
   cos[27]  =  16'b0011111100011111;     //27pi/512
   sin[28]  =  16'b1111010100001111;     //28pi/512
   cos[28]  =  16'b0011111100001110;     //28pi/512
   sin[29]  =  16'b1111010010101100;     //29pi/512
   cos[29]  =  16'b0011111011111101;     //29pi/512
   sin[30]  =  16'b1111010001001001;     //30pi/512
   cos[30]  =  16'b0011111011101011;     //30pi/512
   sin[31]  =  16'b1111001111100110;     //31pi/512
   cos[31]  =  16'b0011111011011000;     //31pi/512
   sin[32]  =  16'b1111001110000100;     //32pi/512
   cos[32]  =  16'b0011111011000101;     //32pi/512
   sin[33]  =  16'b1111001100100001;     //33pi/512
   cos[33]  =  16'b0011111010110001;     //33pi/512
   sin[34]  =  16'b1111001010111111;     //34pi/512
   cos[34]  =  16'b0011111010011100;     //34pi/512
   sin[35]  =  16'b1111001001011100;     //35pi/512
   cos[35]  =  16'b0011111010000111;     //35pi/512
   sin[36]  =  16'b1111000111111010;     //36pi/512
   cos[36]  =  16'b0011111001110001;     //36pi/512
   sin[37]  =  16'b1111000110011000;     //37pi/512
   cos[37]  =  16'b0011111001011011;     //37pi/512
   sin[38]  =  16'b1111000100110110;     //38pi/512
   cos[38]  =  16'b0011111001000100;     //38pi/512
   sin[39]  =  16'b1111000011010101;     //39pi/512
   cos[39]  =  16'b0011111000101101;     //39pi/512
   sin[40]  =  16'b1111000001110011;     //40pi/512
   cos[40]  =  16'b0011111000010100;     //40pi/512
   sin[41]  =  16'b1111000000010010;     //41pi/512
   cos[41]  =  16'b0011110111111100;     //41pi/512
   sin[42]  =  16'b1110111110110000;     //42pi/512
   cos[42]  =  16'b0011110111100010;     //42pi/512
   sin[43]  =  16'b1110111101001111;     //43pi/512
   cos[43]  =  16'b0011110111001001;     //43pi/512
   sin[44]  =  16'b1110111011101110;     //44pi/512
   cos[44]  =  16'b0011110110101110;     //44pi/512
   sin[45]  =  16'b1110111010001101;     //45pi/512
   cos[45]  =  16'b0011110110010011;     //45pi/512
   sin[46]  =  16'b1110111000101101;     //46pi/512
   cos[46]  =  16'b0011110101110111;     //46pi/512
   sin[47]  =  16'b1110110111001100;     //47pi/512
   cos[47]  =  16'b0011110101011011;     //47pi/512
   sin[48]  =  16'b1110110101101100;     //48pi/512
   cos[48]  =  16'b0011110100111110;     //48pi/512
   sin[49]  =  16'b1110110100001100;     //49pi/512
   cos[49]  =  16'b0011110100100001;     //49pi/512
   sin[50]  =  16'b1110110010101100;     //50pi/512
   cos[50]  =  16'b0011110100000010;     //50pi/512
   sin[51]  =  16'b1110110001001100;     //51pi/512
   cos[51]  =  16'b0011110011100100;     //51pi/512
   sin[52]  =  16'b1110101111101101;     //52pi/512
   cos[52]  =  16'b0011110011000101;     //52pi/512
   sin[53]  =  16'b1110101110001101;     //53pi/512
   cos[53]  =  16'b0011110010100101;     //53pi/512
   sin[54]  =  16'b1110101100101110;     //54pi/512
   cos[54]  =  16'b0011110010000100;     //54pi/512
   sin[55]  =  16'b1110101011001111;     //55pi/512
   cos[55]  =  16'b0011110001100011;     //55pi/512
   sin[56]  =  16'b1110101001110000;     //56pi/512
   cos[56]  =  16'b0011110001000010;     //56pi/512
   sin[57]  =  16'b1110101000010010;     //57pi/512
   cos[57]  =  16'b0011110000100000;     //57pi/512
   sin[58]  =  16'b1110100110110100;     //58pi/512
   cos[58]  =  16'b0011101111111101;     //58pi/512
   sin[59]  =  16'b1110100101010101;     //59pi/512
   cos[59]  =  16'b0011101111011010;     //59pi/512
   sin[60]  =  16'b1110100011110111;     //60pi/512
   cos[60]  =  16'b0011101110110110;     //60pi/512
   sin[61]  =  16'b1110100010011010;     //61pi/512
   cos[61]  =  16'b0011101110010001;     //61pi/512
   sin[62]  =  16'b1110100000111100;     //62pi/512
   cos[62]  =  16'b0011101101101100;     //62pi/512
   sin[63]  =  16'b1110011111011111;     //63pi/512
   cos[63]  =  16'b0011101101000111;     //63pi/512
   sin[64]  =  16'b1110011110000010;     //64pi/512
   cos[64]  =  16'b0011101100100000;     //64pi/512
   sin[65]  =  16'b1110011100100101;     //65pi/512
   cos[65]  =  16'b0011101011111010;     //65pi/512
   sin[66]  =  16'b1110011011001001;     //66pi/512
   cos[66]  =  16'b0011101011010010;     //66pi/512
   sin[67]  =  16'b1110011001101101;     //67pi/512
   cos[67]  =  16'b0011101010101010;     //67pi/512
   sin[68]  =  16'b1110011000010001;     //68pi/512
   cos[68]  =  16'b0011101010000010;     //68pi/512
   sin[69]  =  16'b1110010110110101;     //69pi/512
   cos[69]  =  16'b0011101001011001;     //69pi/512
   sin[70]  =  16'b1110010101011001;     //70pi/512
   cos[70]  =  16'b0011101000101111;     //70pi/512
   sin[71]  =  16'b1110010011111110;     //71pi/512
   cos[71]  =  16'b0011101000000101;     //71pi/512
   sin[72]  =  16'b1110010010100011;     //72pi/512
   cos[72]  =  16'b0011100111011010;     //72pi/512
   sin[73]  =  16'b1110010001001000;     //73pi/512
   cos[73]  =  16'b0011100110101111;     //73pi/512
   sin[74]  =  16'b1110001111101110;     //74pi/512
   cos[74]  =  16'b0011100110000011;     //74pi/512
   sin[75]  =  16'b1110001110010100;     //75pi/512
   cos[75]  =  16'b0011100101010111;     //75pi/512
   sin[76]  =  16'b1110001100111010;     //76pi/512
   cos[76]  =  16'b0011100100101010;     //76pi/512
   sin[77]  =  16'b1110001011100000;     //77pi/512
   cos[77]  =  16'b0011100011111101;     //77pi/512
   sin[78]  =  16'b1110001010000111;     //78pi/512
   cos[78]  =  16'b0011100011001111;     //78pi/512
   sin[79]  =  16'b1110001000101101;     //79pi/512
   cos[79]  =  16'b0011100010100000;     //79pi/512
   sin[80]  =  16'b1110000111010101;     //80pi/512
   cos[80]  =  16'b0011100001110001;     //80pi/512
   sin[81]  =  16'b1110000101111100;     //81pi/512
   cos[81]  =  16'b0011100001000001;     //81pi/512
   sin[82]  =  16'b1110000100100100;     //82pi/512
   cos[82]  =  16'b0011100000010001;     //82pi/512
   sin[83]  =  16'b1110000011001100;     //83pi/512
   cos[83]  =  16'b0011011111100000;     //83pi/512
   sin[84]  =  16'b1110000001110100;     //84pi/512
   cos[84]  =  16'b0011011110101111;     //84pi/512
   sin[85]  =  16'b1110000000011101;     //85pi/512
   cos[85]  =  16'b0011011101111101;     //85pi/512
   sin[86]  =  16'b1101111111000110;     //86pi/512
   cos[86]  =  16'b0011011101001011;     //86pi/512
   sin[87]  =  16'b1101111101101111;     //87pi/512
   cos[87]  =  16'b0011011100011000;     //87pi/512
   sin[88]  =  16'b1101111100011001;     //88pi/512
   cos[88]  =  16'b0011011011100101;     //88pi/512
   sin[89]  =  16'b1101111011000011;     //89pi/512
   cos[89]  =  16'b0011011010110001;     //89pi/512
   sin[90]  =  16'b1101111001101101;     //90pi/512
   cos[90]  =  16'b0011011001111100;     //90pi/512
   sin[91]  =  16'b1101111000011000;     //91pi/512
   cos[91]  =  16'b0011011001000111;     //91pi/512
   sin[92]  =  16'b1101110111000011;     //92pi/512
   cos[92]  =  16'b0011011000010010;     //92pi/512
   sin[93]  =  16'b1101110101101110;     //93pi/512
   cos[93]  =  16'b0011010111011100;     //93pi/512
   sin[94]  =  16'b1101110100011001;     //94pi/512
   cos[94]  =  16'b0011010110100101;     //94pi/512
   sin[95]  =  16'b1101110011000101;     //95pi/512
   cos[95]  =  16'b0011010101101110;     //95pi/512
   sin[96]  =  16'b1101110001110010;     //96pi/512
   cos[96]  =  16'b0011010100110110;     //96pi/512
   sin[97]  =  16'b1101110000011110;     //97pi/512
   cos[97]  =  16'b0011010011111110;     //97pi/512
   sin[98]  =  16'b1101101111001011;     //98pi/512
   cos[98]  =  16'b0011010011000110;     //98pi/512
   sin[99]  =  16'b1101101101111000;     //99pi/512
   cos[99]  =  16'b0011010010001100;     //99pi/512
   sin[100]  =  16'b1101101100100110;     //100pi/512
   cos[100]  =  16'b0011010001010011;     //100pi/512
   sin[101]  =  16'b1101101011010100;     //101pi/512
   cos[101]  =  16'b0011010000011001;     //101pi/512
   sin[102]  =  16'b1101101010000010;     //102pi/512
   cos[102]  =  16'b0011001111011110;     //102pi/512
   sin[103]  =  16'b1101101000110001;     //103pi/512
   cos[103]  =  16'b0011001110100011;     //103pi/512
   sin[104]  =  16'b1101100111100000;     //104pi/512
   cos[104]  =  16'b0011001101100111;     //104pi/512
   sin[105]  =  16'b1101100110001111;     //105pi/512
   cos[105]  =  16'b0011001100101011;     //105pi/512
   sin[106]  =  16'b1101100100111111;     //106pi/512
   cos[106]  =  16'b0011001011101110;     //106pi/512
   sin[107]  =  16'b1101100011101111;     //107pi/512
   cos[107]  =  16'b0011001010110001;     //107pi/512
   sin[108]  =  16'b1101100010100000;     //108pi/512
   cos[108]  =  16'b0011001001110100;     //108pi/512
   sin[109]  =  16'b1101100001010001;     //109pi/512
   cos[109]  =  16'b0011001000110110;     //109pi/512
   sin[110]  =  16'b1101100000000010;     //110pi/512
   cos[110]  =  16'b0011000111110111;     //110pi/512
   sin[111]  =  16'b1101011110110100;     //111pi/512
   cos[111]  =  16'b0011000110111000;     //111pi/512
   sin[112]  =  16'b1101011101100110;     //112pi/512
   cos[112]  =  16'b0011000101111001;     //112pi/512
   sin[113]  =  16'b1101011100011001;     //113pi/512
   cos[113]  =  16'b0011000100111000;     //113pi/512
   sin[114]  =  16'b1101011011001011;     //114pi/512
   cos[114]  =  16'b0011000011111000;     //114pi/512
   sin[115]  =  16'b1101011001111111;     //115pi/512
   cos[115]  =  16'b0011000010110111;     //115pi/512
   sin[116]  =  16'b1101011000110010;     //116pi/512
   cos[116]  =  16'b0011000001110110;     //116pi/512
   sin[117]  =  16'b1101010111100110;     //117pi/512
   cos[117]  =  16'b0011000000110100;     //117pi/512
   sin[118]  =  16'b1101010110011011;     //118pi/512
   cos[118]  =  16'b0010111111110001;     //118pi/512
   sin[119]  =  16'b1101010101010000;     //119pi/512
   cos[119]  =  16'b0010111110101111;     //119pi/512
   sin[120]  =  16'b1101010100000101;     //120pi/512
   cos[120]  =  16'b0010111101101011;     //120pi/512
   sin[121]  =  16'b1101010010111011;     //121pi/512
   cos[121]  =  16'b0010111100101000;     //121pi/512
   sin[122]  =  16'b1101010001110001;     //122pi/512
   cos[122]  =  16'b0010111011100011;     //122pi/512
   sin[123]  =  16'b1101010000101000;     //123pi/512
   cos[123]  =  16'b0010111010011111;     //123pi/512
   sin[124]  =  16'b1101001111011111;     //124pi/512
   cos[124]  =  16'b0010111001011010;     //124pi/512
   sin[125]  =  16'b1101001110010110;     //125pi/512
   cos[125]  =  16'b0010111000010100;     //125pi/512
   sin[126]  =  16'b1101001101001110;     //126pi/512
   cos[126]  =  16'b0010110111001110;     //126pi/512
   sin[127]  =  16'b1101001100000110;     //127pi/512
   cos[127]  =  16'b0010110110001000;     //127pi/512
   sin[128]  =  16'b1101001010111111;     //128pi/512
   cos[128]  =  16'b0010110101000001;     //128pi/512
   sin[129]  =  16'b1101001001111000;     //129pi/512
   cos[129]  =  16'b0010110011111001;     //129pi/512
   sin[130]  =  16'b1101001000110001;     //130pi/512
   cos[130]  =  16'b0010110010110010;     //130pi/512
   sin[131]  =  16'b1101000111101011;     //131pi/512
   cos[131]  =  16'b0010110001101010;     //131pi/512
   sin[132]  =  16'b1101000110100110;     //132pi/512
   cos[132]  =  16'b0010110000100001;     //132pi/512
   sin[133]  =  16'b1101000101100001;     //133pi/512
   cos[133]  =  16'b0010101111011000;     //133pi/512
   sin[134]  =  16'b1101000100011100;     //134pi/512
   cos[134]  =  16'b0010101110001110;     //134pi/512
   sin[135]  =  16'b1101000011011000;     //135pi/512
   cos[135]  =  16'b0010101101000101;     //135pi/512
   sin[136]  =  16'b1101000010010100;     //136pi/512
   cos[136]  =  16'b0010101011111010;     //136pi/512
   sin[137]  =  16'b1101000001010001;     //137pi/512
   cos[137]  =  16'b0010101010110000;     //137pi/512
   sin[138]  =  16'b1101000000001110;     //138pi/512
   cos[138]  =  16'b0010101001100101;     //138pi/512
   sin[139]  =  16'b1100111111001100;     //139pi/512
   cos[139]  =  16'b0010101000011001;     //139pi/512
   sin[140]  =  16'b1100111110001010;     //140pi/512
   cos[140]  =  16'b0010100111001101;     //140pi/512
   sin[141]  =  16'b1100111101001000;     //141pi/512
   cos[141]  =  16'b0010100110000001;     //141pi/512
   sin[142]  =  16'b1100111100000111;     //142pi/512
   cos[142]  =  16'b0010100100110100;     //142pi/512
   sin[143]  =  16'b1100111011000111;     //143pi/512
   cos[143]  =  16'b0010100011100111;     //143pi/512
   sin[144]  =  16'b1100111010000111;     //144pi/512
   cos[144]  =  16'b0010100010011001;     //144pi/512
   sin[145]  =  16'b1100111001000111;     //145pi/512
   cos[145]  =  16'b0010100001001011;     //145pi/512
   sin[146]  =  16'b1100111000001000;     //146pi/512
   cos[146]  =  16'b0010011111111101;     //146pi/512
   sin[147]  =  16'b1100110111001010;     //147pi/512
   cos[147]  =  16'b0010011110101111;     //147pi/512
   sin[148]  =  16'b1100110110001100;     //148pi/512
   cos[148]  =  16'b0010011101011111;     //148pi/512
   sin[149]  =  16'b1100110101001110;     //149pi/512
   cos[149]  =  16'b0010011100010000;     //149pi/512
   sin[150]  =  16'b1100110100010001;     //150pi/512
   cos[150]  =  16'b0010011011000000;     //150pi/512
   sin[151]  =  16'b1100110011010100;     //151pi/512
   cos[151]  =  16'b0010011001110000;     //151pi/512
   sin[152]  =  16'b1100110010011000;     //152pi/512
   cos[152]  =  16'b0010011000011111;     //152pi/512
   sin[153]  =  16'b1100110001011101;     //153pi/512
   cos[153]  =  16'b0010010111001111;     //153pi/512
   sin[154]  =  16'b1100110000100001;     //154pi/512
   cos[154]  =  16'b0010010101111101;     //154pi/512
   sin[155]  =  16'b1100101111100111;     //155pi/512
   cos[155]  =  16'b0010010100101100;     //155pi/512
   sin[156]  =  16'b1100101110101101;     //156pi/512
   cos[156]  =  16'b0010010011011010;     //156pi/512
   sin[157]  =  16'b1100101101110011;     //157pi/512
   cos[157]  =  16'b0010010010000111;     //157pi/512
   sin[158]  =  16'b1100101100111010;     //158pi/512
   cos[158]  =  16'b0010010000110100;     //158pi/512
   sin[159]  =  16'b1100101100000001;     //159pi/512
   cos[159]  =  16'b0010001111100001;     //159pi/512
   sin[160]  =  16'b1100101011001001;     //160pi/512
   cos[160]  =  16'b0010001110001110;     //160pi/512
   sin[161]  =  16'b1100101010010010;     //161pi/512
   cos[161]  =  16'b0010001100111010;     //161pi/512
   sin[162]  =  16'b1100101001011011;     //162pi/512
   cos[162]  =  16'b0010001011100110;     //162pi/512
   sin[163]  =  16'b1100101000100100;     //163pi/512
   cos[163]  =  16'b0010001010010010;     //163pi/512
   sin[164]  =  16'b1100100111101110;     //164pi/512
   cos[164]  =  16'b0010001000111101;     //164pi/512
   sin[165]  =  16'b1100100110111000;     //165pi/512
   cos[165]  =  16'b0010000111101000;     //165pi/512
   sin[166]  =  16'b1100100110000011;     //166pi/512
   cos[166]  =  16'b0010000110010010;     //166pi/512
   sin[167]  =  16'b1100100101001111;     //167pi/512
   cos[167]  =  16'b0010000100111101;     //167pi/512
   sin[168]  =  16'b1100100100011011;     //168pi/512
   cos[168]  =  16'b0010000011100111;     //168pi/512
   sin[169]  =  16'b1100100011101000;     //169pi/512
   cos[169]  =  16'b0010000010010000;     //169pi/512
   sin[170]  =  16'b1100100010110101;     //170pi/512
   cos[170]  =  16'b0010000000111001;     //170pi/512
   sin[171]  =  16'b1100100010000010;     //171pi/512
   cos[171]  =  16'b0001111111100010;     //171pi/512
   sin[172]  =  16'b1100100001010000;     //172pi/512
   cos[172]  =  16'b0001111110001011;     //172pi/512
   sin[173]  =  16'b1100100000011111;     //173pi/512
   cos[173]  =  16'b0001111100110100;     //173pi/512
   sin[174]  =  16'b1100011111101110;     //174pi/512
   cos[174]  =  16'b0001111011011100;     //174pi/512
   sin[175]  =  16'b1100011110111110;     //175pi/512
   cos[175]  =  16'b0001111010000011;     //175pi/512
   sin[176]  =  16'b1100011110001111;     //176pi/512
   cos[176]  =  16'b0001111000101011;     //176pi/512
   sin[177]  =  16'b1100011101011111;     //177pi/512
   cos[177]  =  16'b0001110111010010;     //177pi/512
   sin[178]  =  16'b1100011100110001;     //178pi/512
   cos[178]  =  16'b0001110101111001;     //178pi/512
   sin[179]  =  16'b1100011100000011;     //179pi/512
   cos[179]  =  16'b0001110100100000;     //179pi/512
   sin[180]  =  16'b1100011011010101;     //180pi/512
   cos[180]  =  16'b0001110011000110;     //180pi/512
   sin[181]  =  16'b1100011010101000;     //181pi/512
   cos[181]  =  16'b0001110001101100;     //181pi/512
   sin[182]  =  16'b1100011001111100;     //182pi/512
   cos[182]  =  16'b0001110000010010;     //182pi/512
   sin[183]  =  16'b1100011001010000;     //183pi/512
   cos[183]  =  16'b0001101110110111;     //183pi/512
   sin[184]  =  16'b1100011000100101;     //184pi/512
   cos[184]  =  16'b0001101101011101;     //184pi/512
   sin[185]  =  16'b1100010111111010;     //185pi/512
   cos[185]  =  16'b0001101100000010;     //185pi/512
   sin[186]  =  16'b1100010111010000;     //186pi/512
   cos[186]  =  16'b0001101010100110;     //186pi/512
   sin[187]  =  16'b1100010110100111;     //187pi/512
   cos[187]  =  16'b0001101001001011;     //187pi/512
   sin[188]  =  16'b1100010101111110;     //188pi/512
   cos[188]  =  16'b0001100111101111;     //188pi/512
   sin[189]  =  16'b1100010101010101;     //189pi/512
   cos[189]  =  16'b0001100110010011;     //189pi/512
   sin[190]  =  16'b1100010100101101;     //190pi/512
   cos[190]  =  16'b0001100100110111;     //190pi/512
   sin[191]  =  16'b1100010100000110;     //191pi/512
   cos[191]  =  16'b0001100011011010;     //191pi/512
   sin[192]  =  16'b1100010011011111;     //192pi/512
   cos[192]  =  16'b0001100001111101;     //192pi/512
   sin[193]  =  16'b1100010010111001;     //193pi/512
   cos[193]  =  16'b0001100000100000;     //193pi/512
   sin[194]  =  16'b1100010010010011;     //194pi/512
   cos[194]  =  16'b0001011111000011;     //194pi/512
   sin[195]  =  16'b1100010001101110;     //195pi/512
   cos[195]  =  16'b0001011101100110;     //195pi/512
   sin[196]  =  16'b1100010001001010;     //196pi/512
   cos[196]  =  16'b0001011100001000;     //196pi/512
   sin[197]  =  16'b1100010000100110;     //197pi/512
   cos[197]  =  16'b0001011010101010;     //197pi/512
   sin[198]  =  16'b1100010000000011;     //198pi/512
   cos[198]  =  16'b0001011001001100;     //198pi/512
   sin[199]  =  16'b1100001111100000;     //199pi/512
   cos[199]  =  16'b0001010111101110;     //199pi/512
   sin[200]  =  16'b1100001110111110;     //200pi/512
   cos[200]  =  16'b0001010110001111;     //200pi/512
   sin[201]  =  16'b1100001110011100;     //201pi/512
   cos[201]  =  16'b0001010100110000;     //201pi/512
   sin[202]  =  16'b1100001101111011;     //202pi/512
   cos[202]  =  16'b0001010011010001;     //202pi/512
   sin[203]  =  16'b1100001101011011;     //203pi/512
   cos[203]  =  16'b0001010001110010;     //203pi/512
   sin[204]  =  16'b1100001100111011;     //204pi/512
   cos[204]  =  16'b0001010000010011;     //204pi/512
   sin[205]  =  16'b1100001100011100;     //205pi/512
   cos[205]  =  16'b0001001110110011;     //205pi/512
   sin[206]  =  16'b1100001011111101;     //206pi/512
   cos[206]  =  16'b0001001101010100;     //206pi/512
   sin[207]  =  16'b1100001011011111;     //207pi/512
   cos[207]  =  16'b0001001011110100;     //207pi/512
   sin[208]  =  16'b1100001011000001;     //208pi/512
   cos[208]  =  16'b0001001010010100;     //208pi/512
   sin[209]  =  16'b1100001010100101;     //209pi/512
   cos[209]  =  16'b0001001000110011;     //209pi/512
   sin[210]  =  16'b1100001010001000;     //210pi/512
   cos[210]  =  16'b0001000111010011;     //210pi/512
   sin[211]  =  16'b1100001001101101;     //211pi/512
   cos[211]  =  16'b0001000101110010;     //211pi/512
   sin[212]  =  16'b1100001001010001;     //212pi/512
   cos[212]  =  16'b0001000100010001;     //212pi/512
   sin[213]  =  16'b1100001000110111;     //213pi/512
   cos[213]  =  16'b0001000010110000;     //213pi/512
   sin[214]  =  16'b1100001000011101;     //214pi/512
   cos[214]  =  16'b0001000001001111;     //214pi/512
   sin[215]  =  16'b1100001000000100;     //215pi/512
   cos[215]  =  16'b0000111111101110;     //215pi/512
   sin[216]  =  16'b1100000111101011;     //216pi/512
   cos[216]  =  16'b0000111110001100;     //216pi/512
   sin[217]  =  16'b1100000111010011;     //217pi/512
   cos[217]  =  16'b0000111100101011;     //217pi/512
   sin[218]  =  16'b1100000110111011;     //218pi/512
   cos[218]  =  16'b0000111011001001;     //218pi/512
   sin[219]  =  16'b1100000110100100;     //219pi/512
   cos[219]  =  16'b0000111001100111;     //219pi/512
   sin[220]  =  16'b1100000110001110;     //220pi/512
   cos[220]  =  16'b0000111000000101;     //220pi/512
   sin[221]  =  16'b1100000101111000;     //221pi/512
   cos[221]  =  16'b0000110110100011;     //221pi/512
   sin[222]  =  16'b1100000101100011;     //222pi/512
   cos[222]  =  16'b0000110101000001;     //222pi/512
   sin[223]  =  16'b1100000101001111;     //223pi/512
   cos[223]  =  16'b0000110011011110;     //223pi/512
   sin[224]  =  16'b1100000100111011;     //224pi/512
   cos[224]  =  16'b0000110001111100;     //224pi/512
   sin[225]  =  16'b1100000100101000;     //225pi/512
   cos[225]  =  16'b0000110000011001;     //225pi/512
   sin[226]  =  16'b1100000100010101;     //226pi/512
   cos[226]  =  16'b0000101110110110;     //226pi/512
   sin[227]  =  16'b1100000100000011;     //227pi/512
   cos[227]  =  16'b0000101101010100;     //227pi/512
   sin[228]  =  16'b1100000011110001;     //228pi/512
   cos[228]  =  16'b0000101011110001;     //228pi/512
   sin[229]  =  16'b1100000011100000;     //229pi/512
   cos[229]  =  16'b0000101010001101;     //229pi/512
   sin[230]  =  16'b1100000011010000;     //230pi/512
   cos[230]  =  16'b0000101000101010;     //230pi/512
   sin[231]  =  16'b1100000011000000;     //231pi/512
   cos[231]  =  16'b0000100111000111;     //231pi/512
   sin[232]  =  16'b1100000010110001;     //232pi/512
   cos[232]  =  16'b0000100101100100;     //232pi/512
   sin[233]  =  16'b1100000010100011;     //233pi/512
   cos[233]  =  16'b0000100100000000;     //233pi/512
   sin[234]  =  16'b1100000010010101;     //234pi/512
   cos[234]  =  16'b0000100010011100;     //234pi/512
   sin[235]  =  16'b1100000010001000;     //235pi/512
   cos[235]  =  16'b0000100000111001;     //235pi/512
   sin[236]  =  16'b1100000001111011;     //236pi/512
   cos[236]  =  16'b0000011111010101;     //236pi/512
   sin[237]  =  16'b1100000001101111;     //237pi/512
   cos[237]  =  16'b0000011101110001;     //237pi/512
   sin[238]  =  16'b1100000001100100;     //238pi/512
   cos[238]  =  16'b0000011100001101;     //238pi/512
   sin[239]  =  16'b1100000001011001;     //239pi/512
   cos[239]  =  16'b0000011010101001;     //239pi/512
   sin[240]  =  16'b1100000001001111;     //240pi/512
   cos[240]  =  16'b0000011001000101;     //240pi/512
   sin[241]  =  16'b1100000001000101;     //241pi/512
   cos[241]  =  16'b0000010111100001;     //241pi/512
   sin[242]  =  16'b1100000000111100;     //242pi/512
   cos[242]  =  16'b0000010101111101;     //242pi/512
   sin[243]  =  16'b1100000000110100;     //243pi/512
   cos[243]  =  16'b0000010100011001;     //243pi/512
   sin[244]  =  16'b1100000000101100;     //244pi/512
   cos[244]  =  16'b0000010010110101;     //244pi/512
   sin[245]  =  16'b1100000000100101;     //245pi/512
   cos[245]  =  16'b0000010001010001;     //245pi/512
   sin[246]  =  16'b1100000000011111;     //246pi/512
   cos[246]  =  16'b0000001111101100;     //246pi/512
   sin[247]  =  16'b1100000000011001;     //247pi/512
   cos[247]  =  16'b0000001110001000;     //247pi/512
   sin[248]  =  16'b1100000000010100;     //248pi/512
   cos[248]  =  16'b0000001100100011;     //248pi/512
   sin[249]  =  16'b1100000000001111;     //249pi/512
   cos[249]  =  16'b0000001010111111;     //249pi/512
   sin[250]  =  16'b1100000000001011;     //250pi/512
   cos[250]  =  16'b0000001001011011;     //250pi/512
   sin[251]  =  16'b1100000000001000;     //251pi/512
   cos[251]  =  16'b0000000111110110;     //251pi/512
   sin[252]  =  16'b1100000000000101;     //252pi/512
   cos[252]  =  16'b0000000110010010;     //252pi/512
   sin[253]  =  16'b1100000000000011;     //253pi/512
   cos[253]  =  16'b0000000100101101;     //253pi/512
   sin[254]  =  16'b1100000000000001;     //254pi/512
   cos[254]  =  16'b0000000011001001;     //254pi/512
   sin[255]  =  16'b1100000000000000;     //255pi/512
   cos[255]  =  16'b0000000001100100;     //255pi/512
   sin[256]  =  16'b1100000000000000;     //256pi/512
   cos[256]  =  16'b0000000000000000;     //256pi/512
   sin[257]  =  16'b1100000000000000;     //257pi/512
   cos[257]  =  16'b1111111110011011;     //257pi/512
   sin[258]  =  16'b1100000000000001;     //258pi/512
   cos[258]  =  16'b1111111100110111;     //258pi/512
   sin[259]  =  16'b1100000000000011;     //259pi/512
   cos[259]  =  16'b1111111011010010;     //259pi/512
   sin[260]  =  16'b1100000000000101;     //260pi/512
   cos[260]  =  16'b1111111001101110;     //260pi/512
   sin[261]  =  16'b1100000000001000;     //261pi/512
   cos[261]  =  16'b1111111000001001;     //261pi/512
   sin[262]  =  16'b1100000000001011;     //262pi/512
   cos[262]  =  16'b1111110110100101;     //262pi/512
   sin[263]  =  16'b1100000000001111;     //263pi/512
   cos[263]  =  16'b1111110101000000;     //263pi/512
   sin[264]  =  16'b1100000000010100;     //264pi/512
   cos[264]  =  16'b1111110011011100;     //264pi/512
   sin[265]  =  16'b1100000000011001;     //265pi/512
   cos[265]  =  16'b1111110001111000;     //265pi/512
   sin[266]  =  16'b1100000000011111;     //266pi/512
   cos[266]  =  16'b1111110000010011;     //266pi/512
   sin[267]  =  16'b1100000000100101;     //267pi/512
   cos[267]  =  16'b1111101110101111;     //267pi/512
   sin[268]  =  16'b1100000000101100;     //268pi/512
   cos[268]  =  16'b1111101101001011;     //268pi/512
   sin[269]  =  16'b1100000000110100;     //269pi/512
   cos[269]  =  16'b1111101011100110;     //269pi/512
   sin[270]  =  16'b1100000000111100;     //270pi/512
   cos[270]  =  16'b1111101010000010;     //270pi/512
   sin[271]  =  16'b1100000001000101;     //271pi/512
   cos[271]  =  16'b1111101000011110;     //271pi/512
   sin[272]  =  16'b1100000001001111;     //272pi/512
   cos[272]  =  16'b1111100110111010;     //272pi/512
   sin[273]  =  16'b1100000001011001;     //273pi/512
   cos[273]  =  16'b1111100101010110;     //273pi/512
   sin[274]  =  16'b1100000001100100;     //274pi/512
   cos[274]  =  16'b1111100011110010;     //274pi/512
   sin[275]  =  16'b1100000001101111;     //275pi/512
   cos[275]  =  16'b1111100010001110;     //275pi/512
   sin[276]  =  16'b1100000001111011;     //276pi/512
   cos[276]  =  16'b1111100000101010;     //276pi/512
   sin[277]  =  16'b1100000010001000;     //277pi/512
   cos[277]  =  16'b1111011111000111;     //277pi/512
   sin[278]  =  16'b1100000010010101;     //278pi/512
   cos[278]  =  16'b1111011101100011;     //278pi/512
   sin[279]  =  16'b1100000010100011;     //279pi/512
   cos[279]  =  16'b1111011011111111;     //279pi/512
   sin[280]  =  16'b1100000010110001;     //280pi/512
   cos[280]  =  16'b1111011010011100;     //280pi/512
   sin[281]  =  16'b1100000011000000;     //281pi/512
   cos[281]  =  16'b1111011000111001;     //281pi/512
   sin[282]  =  16'b1100000011010000;     //282pi/512
   cos[282]  =  16'b1111010111010101;     //282pi/512
   sin[283]  =  16'b1100000011100000;     //283pi/512
   cos[283]  =  16'b1111010101110010;     //283pi/512
   sin[284]  =  16'b1100000011110001;     //284pi/512
   cos[284]  =  16'b1111010100001111;     //284pi/512
   sin[285]  =  16'b1100000100000011;     //285pi/512
   cos[285]  =  16'b1111010010101100;     //285pi/512
   sin[286]  =  16'b1100000100010101;     //286pi/512
   cos[286]  =  16'b1111010001001001;     //286pi/512
   sin[287]  =  16'b1100000100101000;     //287pi/512
   cos[287]  =  16'b1111001111100110;     //287pi/512
   sin[288]  =  16'b1100000100111011;     //288pi/512
   cos[288]  =  16'b1111001110000100;     //288pi/512
   sin[289]  =  16'b1100000101001111;     //289pi/512
   cos[289]  =  16'b1111001100100001;     //289pi/512
   sin[290]  =  16'b1100000101100011;     //290pi/512
   cos[290]  =  16'b1111001010111111;     //290pi/512
   sin[291]  =  16'b1100000101111000;     //291pi/512
   cos[291]  =  16'b1111001001011100;     //291pi/512
   sin[292]  =  16'b1100000110001110;     //292pi/512
   cos[292]  =  16'b1111000111111010;     //292pi/512
   sin[293]  =  16'b1100000110100100;     //293pi/512
   cos[293]  =  16'b1111000110011000;     //293pi/512
   sin[294]  =  16'b1100000110111011;     //294pi/512
   cos[294]  =  16'b1111000100110110;     //294pi/512
   sin[295]  =  16'b1100000111010011;     //295pi/512
   cos[295]  =  16'b1111000011010101;     //295pi/512
   sin[296]  =  16'b1100000111101011;     //296pi/512
   cos[296]  =  16'b1111000001110011;     //296pi/512
   sin[297]  =  16'b1100001000000100;     //297pi/512
   cos[297]  =  16'b1111000000010010;     //297pi/512
   sin[298]  =  16'b1100001000011101;     //298pi/512
   cos[298]  =  16'b1110111110110000;     //298pi/512
   sin[299]  =  16'b1100001000110111;     //299pi/512
   cos[299]  =  16'b1110111101001111;     //299pi/512
   sin[300]  =  16'b1100001001010001;     //300pi/512
   cos[300]  =  16'b1110111011101110;     //300pi/512
   sin[301]  =  16'b1100001001101101;     //301pi/512
   cos[301]  =  16'b1110111010001101;     //301pi/512
   sin[302]  =  16'b1100001010001000;     //302pi/512
   cos[302]  =  16'b1110111000101101;     //302pi/512
   sin[303]  =  16'b1100001010100101;     //303pi/512
   cos[303]  =  16'b1110110111001100;     //303pi/512
   sin[304]  =  16'b1100001011000001;     //304pi/512
   cos[304]  =  16'b1110110101101100;     //304pi/512
   sin[305]  =  16'b1100001011011111;     //305pi/512
   cos[305]  =  16'b1110110100001100;     //305pi/512
   sin[306]  =  16'b1100001011111101;     //306pi/512
   cos[306]  =  16'b1110110010101100;     //306pi/512
   sin[307]  =  16'b1100001100011100;     //307pi/512
   cos[307]  =  16'b1110110001001100;     //307pi/512
   sin[308]  =  16'b1100001100111011;     //308pi/512
   cos[308]  =  16'b1110101111101101;     //308pi/512
   sin[309]  =  16'b1100001101011011;     //309pi/512
   cos[309]  =  16'b1110101110001101;     //309pi/512
   sin[310]  =  16'b1100001101111011;     //310pi/512
   cos[310]  =  16'b1110101100101110;     //310pi/512
   sin[311]  =  16'b1100001110011100;     //311pi/512
   cos[311]  =  16'b1110101011001111;     //311pi/512
   sin[312]  =  16'b1100001110111110;     //312pi/512
   cos[312]  =  16'b1110101001110000;     //312pi/512
   sin[313]  =  16'b1100001111100000;     //313pi/512
   cos[313]  =  16'b1110101000010010;     //313pi/512
   sin[314]  =  16'b1100010000000011;     //314pi/512
   cos[314]  =  16'b1110100110110100;     //314pi/512
   sin[315]  =  16'b1100010000100110;     //315pi/512
   cos[315]  =  16'b1110100101010101;     //315pi/512
   sin[316]  =  16'b1100010001001010;     //316pi/512
   cos[316]  =  16'b1110100011110111;     //316pi/512
   sin[317]  =  16'b1100010001101110;     //317pi/512
   cos[317]  =  16'b1110100010011010;     //317pi/512
   sin[318]  =  16'b1100010010010011;     //318pi/512
   cos[318]  =  16'b1110100000111100;     //318pi/512
   sin[319]  =  16'b1100010010111001;     //319pi/512
   cos[319]  =  16'b1110011111011111;     //319pi/512
   sin[320]  =  16'b1100010011011111;     //320pi/512
   cos[320]  =  16'b1110011110000010;     //320pi/512
   sin[321]  =  16'b1100010100000110;     //321pi/512
   cos[321]  =  16'b1110011100100101;     //321pi/512
   sin[322]  =  16'b1100010100101101;     //322pi/512
   cos[322]  =  16'b1110011011001001;     //322pi/512
   sin[323]  =  16'b1100010101010101;     //323pi/512
   cos[323]  =  16'b1110011001101101;     //323pi/512
   sin[324]  =  16'b1100010101111110;     //324pi/512
   cos[324]  =  16'b1110011000010001;     //324pi/512
   sin[325]  =  16'b1100010110100111;     //325pi/512
   cos[325]  =  16'b1110010110110101;     //325pi/512
   sin[326]  =  16'b1100010111010000;     //326pi/512
   cos[326]  =  16'b1110010101011001;     //326pi/512
   sin[327]  =  16'b1100010111111010;     //327pi/512
   cos[327]  =  16'b1110010011111110;     //327pi/512
   sin[328]  =  16'b1100011000100101;     //328pi/512
   cos[328]  =  16'b1110010010100011;     //328pi/512
   sin[329]  =  16'b1100011001010000;     //329pi/512
   cos[329]  =  16'b1110010001001000;     //329pi/512
   sin[330]  =  16'b1100011001111100;     //330pi/512
   cos[330]  =  16'b1110001111101110;     //330pi/512
   sin[331]  =  16'b1100011010101000;     //331pi/512
   cos[331]  =  16'b1110001110010100;     //331pi/512
   sin[332]  =  16'b1100011011010101;     //332pi/512
   cos[332]  =  16'b1110001100111010;     //332pi/512
   sin[333]  =  16'b1100011100000011;     //333pi/512
   cos[333]  =  16'b1110001011100000;     //333pi/512
   sin[334]  =  16'b1100011100110001;     //334pi/512
   cos[334]  =  16'b1110001010000111;     //334pi/512
   sin[335]  =  16'b1100011101011111;     //335pi/512
   cos[335]  =  16'b1110001000101101;     //335pi/512
   sin[336]  =  16'b1100011110001111;     //336pi/512
   cos[336]  =  16'b1110000111010101;     //336pi/512
   sin[337]  =  16'b1100011110111110;     //337pi/512
   cos[337]  =  16'b1110000101111100;     //337pi/512
   sin[338]  =  16'b1100011111101110;     //338pi/512
   cos[338]  =  16'b1110000100100100;     //338pi/512
   sin[339]  =  16'b1100100000011111;     //339pi/512
   cos[339]  =  16'b1110000011001100;     //339pi/512
   sin[340]  =  16'b1100100001010000;     //340pi/512
   cos[340]  =  16'b1110000001110100;     //340pi/512
   sin[341]  =  16'b1100100010000010;     //341pi/512
   cos[341]  =  16'b1110000000011101;     //341pi/512
   sin[342]  =  16'b1100100010110101;     //342pi/512
   cos[342]  =  16'b1101111111000110;     //342pi/512
   sin[343]  =  16'b1100100011101000;     //343pi/512
   cos[343]  =  16'b1101111101101111;     //343pi/512
   sin[344]  =  16'b1100100100011011;     //344pi/512
   cos[344]  =  16'b1101111100011001;     //344pi/512
   sin[345]  =  16'b1100100101001111;     //345pi/512
   cos[345]  =  16'b1101111011000011;     //345pi/512
   sin[346]  =  16'b1100100110000011;     //346pi/512
   cos[346]  =  16'b1101111001101101;     //346pi/512
   sin[347]  =  16'b1100100110111000;     //347pi/512
   cos[347]  =  16'b1101111000011000;     //347pi/512
   sin[348]  =  16'b1100100111101110;     //348pi/512
   cos[348]  =  16'b1101110111000011;     //348pi/512
   sin[349]  =  16'b1100101000100100;     //349pi/512
   cos[349]  =  16'b1101110101101110;     //349pi/512
   sin[350]  =  16'b1100101001011011;     //350pi/512
   cos[350]  =  16'b1101110100011001;     //350pi/512
   sin[351]  =  16'b1100101010010010;     //351pi/512
   cos[351]  =  16'b1101110011000101;     //351pi/512
   sin[352]  =  16'b1100101011001001;     //352pi/512
   cos[352]  =  16'b1101110001110010;     //352pi/512
   sin[353]  =  16'b1100101100000001;     //353pi/512
   cos[353]  =  16'b1101110000011110;     //353pi/512
   sin[354]  =  16'b1100101100111010;     //354pi/512
   cos[354]  =  16'b1101101111001011;     //354pi/512
   sin[355]  =  16'b1100101101110011;     //355pi/512
   cos[355]  =  16'b1101101101111000;     //355pi/512
   sin[356]  =  16'b1100101110101101;     //356pi/512
   cos[356]  =  16'b1101101100100110;     //356pi/512
   sin[357]  =  16'b1100101111100111;     //357pi/512
   cos[357]  =  16'b1101101011010100;     //357pi/512
   sin[358]  =  16'b1100110000100001;     //358pi/512
   cos[358]  =  16'b1101101010000010;     //358pi/512
   sin[359]  =  16'b1100110001011101;     //359pi/512
   cos[359]  =  16'b1101101000110001;     //359pi/512
   sin[360]  =  16'b1100110010011000;     //360pi/512
   cos[360]  =  16'b1101100111100000;     //360pi/512
   sin[361]  =  16'b1100110011010100;     //361pi/512
   cos[361]  =  16'b1101100110001111;     //361pi/512
   sin[362]  =  16'b1100110100010001;     //362pi/512
   cos[362]  =  16'b1101100100111111;     //362pi/512
   sin[363]  =  16'b1100110101001110;     //363pi/512
   cos[363]  =  16'b1101100011101111;     //363pi/512
   sin[364]  =  16'b1100110110001100;     //364pi/512
   cos[364]  =  16'b1101100010100000;     //364pi/512
   sin[365]  =  16'b1100110111001010;     //365pi/512
   cos[365]  =  16'b1101100001010001;     //365pi/512
   sin[366]  =  16'b1100111000001000;     //366pi/512
   cos[366]  =  16'b1101100000000010;     //366pi/512
   sin[367]  =  16'b1100111001000111;     //367pi/512
   cos[367]  =  16'b1101011110110100;     //367pi/512
   sin[368]  =  16'b1100111010000111;     //368pi/512
   cos[368]  =  16'b1101011101100110;     //368pi/512
   sin[369]  =  16'b1100111011000111;     //369pi/512
   cos[369]  =  16'b1101011100011001;     //369pi/512
   sin[370]  =  16'b1100111100000111;     //370pi/512
   cos[370]  =  16'b1101011011001011;     //370pi/512
   sin[371]  =  16'b1100111101001000;     //371pi/512
   cos[371]  =  16'b1101011001111111;     //371pi/512
   sin[372]  =  16'b1100111110001010;     //372pi/512
   cos[372]  =  16'b1101011000110010;     //372pi/512
   sin[373]  =  16'b1100111111001100;     //373pi/512
   cos[373]  =  16'b1101010111100110;     //373pi/512
   sin[374]  =  16'b1101000000001110;     //374pi/512
   cos[374]  =  16'b1101010110011011;     //374pi/512
   sin[375]  =  16'b1101000001010001;     //375pi/512
   cos[375]  =  16'b1101010101010000;     //375pi/512
   sin[376]  =  16'b1101000010010100;     //376pi/512
   cos[376]  =  16'b1101010100000101;     //376pi/512
   sin[377]  =  16'b1101000011011000;     //377pi/512
   cos[377]  =  16'b1101010010111011;     //377pi/512
   sin[378]  =  16'b1101000100011100;     //378pi/512
   cos[378]  =  16'b1101010001110001;     //378pi/512
   sin[379]  =  16'b1101000101100001;     //379pi/512
   cos[379]  =  16'b1101010000101000;     //379pi/512
   sin[380]  =  16'b1101000110100110;     //380pi/512
   cos[380]  =  16'b1101001111011111;     //380pi/512
   sin[381]  =  16'b1101000111101011;     //381pi/512
   cos[381]  =  16'b1101001110010110;     //381pi/512
   sin[382]  =  16'b1101001000110001;     //382pi/512
   cos[382]  =  16'b1101001101001110;     //382pi/512
   sin[383]  =  16'b1101001001111000;     //383pi/512
   cos[383]  =  16'b1101001100000110;     //383pi/512
   sin[384]  =  16'b1101001010111111;     //384pi/512
   cos[384]  =  16'b1101001010111111;     //384pi/512
   sin[385]  =  16'b1101001100000110;     //385pi/512
   cos[385]  =  16'b1101001001111000;     //385pi/512
   sin[386]  =  16'b1101001101001110;     //386pi/512
   cos[386]  =  16'b1101001000110001;     //386pi/512
   sin[387]  =  16'b1101001110010110;     //387pi/512
   cos[387]  =  16'b1101000111101011;     //387pi/512
   sin[388]  =  16'b1101001111011111;     //388pi/512
   cos[388]  =  16'b1101000110100110;     //388pi/512
   sin[389]  =  16'b1101010000101000;     //389pi/512
   cos[389]  =  16'b1101000101100001;     //389pi/512
   sin[390]  =  16'b1101010001110001;     //390pi/512
   cos[390]  =  16'b1101000100011100;     //390pi/512
   sin[391]  =  16'b1101010010111011;     //391pi/512
   cos[391]  =  16'b1101000011011000;     //391pi/512
   sin[392]  =  16'b1101010100000101;     //392pi/512
   cos[392]  =  16'b1101000010010100;     //392pi/512
   sin[393]  =  16'b1101010101010000;     //393pi/512
   cos[393]  =  16'b1101000001010001;     //393pi/512
   sin[394]  =  16'b1101010110011011;     //394pi/512
   cos[394]  =  16'b1101000000001110;     //394pi/512
   sin[395]  =  16'b1101010111100110;     //395pi/512
   cos[395]  =  16'b1100111111001100;     //395pi/512
   sin[396]  =  16'b1101011000110010;     //396pi/512
   cos[396]  =  16'b1100111110001010;     //396pi/512
   sin[397]  =  16'b1101011001111111;     //397pi/512
   cos[397]  =  16'b1100111101001000;     //397pi/512
   sin[398]  =  16'b1101011011001011;     //398pi/512
   cos[398]  =  16'b1100111100000111;     //398pi/512
   sin[399]  =  16'b1101011100011001;     //399pi/512
   cos[399]  =  16'b1100111011000111;     //399pi/512
   sin[400]  =  16'b1101011101100110;     //400pi/512
   cos[400]  =  16'b1100111010000111;     //400pi/512
   sin[401]  =  16'b1101011110110100;     //401pi/512
   cos[401]  =  16'b1100111001000111;     //401pi/512
   sin[402]  =  16'b1101100000000010;     //402pi/512
   cos[402]  =  16'b1100111000001000;     //402pi/512
   sin[403]  =  16'b1101100001010001;     //403pi/512
   cos[403]  =  16'b1100110111001010;     //403pi/512
   sin[404]  =  16'b1101100010100000;     //404pi/512
   cos[404]  =  16'b1100110110001100;     //404pi/512
   sin[405]  =  16'b1101100011101111;     //405pi/512
   cos[405]  =  16'b1100110101001110;     //405pi/512
   sin[406]  =  16'b1101100100111111;     //406pi/512
   cos[406]  =  16'b1100110100010001;     //406pi/512
   sin[407]  =  16'b1101100110001111;     //407pi/512
   cos[407]  =  16'b1100110011010100;     //407pi/512
   sin[408]  =  16'b1101100111100000;     //408pi/512
   cos[408]  =  16'b1100110010011000;     //408pi/512
   sin[409]  =  16'b1101101000110001;     //409pi/512
   cos[409]  =  16'b1100110001011101;     //409pi/512
   sin[410]  =  16'b1101101010000010;     //410pi/512
   cos[410]  =  16'b1100110000100001;     //410pi/512
   sin[411]  =  16'b1101101011010100;     //411pi/512
   cos[411]  =  16'b1100101111100111;     //411pi/512
   sin[412]  =  16'b1101101100100110;     //412pi/512
   cos[412]  =  16'b1100101110101101;     //412pi/512
   sin[413]  =  16'b1101101101111000;     //413pi/512
   cos[413]  =  16'b1100101101110011;     //413pi/512
   sin[414]  =  16'b1101101111001011;     //414pi/512
   cos[414]  =  16'b1100101100111010;     //414pi/512
   sin[415]  =  16'b1101110000011110;     //415pi/512
   cos[415]  =  16'b1100101100000001;     //415pi/512
   sin[416]  =  16'b1101110001110010;     //416pi/512
   cos[416]  =  16'b1100101011001001;     //416pi/512
   sin[417]  =  16'b1101110011000101;     //417pi/512
   cos[417]  =  16'b1100101010010010;     //417pi/512
   sin[418]  =  16'b1101110100011001;     //418pi/512
   cos[418]  =  16'b1100101001011011;     //418pi/512
   sin[419]  =  16'b1101110101101110;     //419pi/512
   cos[419]  =  16'b1100101000100100;     //419pi/512
   sin[420]  =  16'b1101110111000011;     //420pi/512
   cos[420]  =  16'b1100100111101110;     //420pi/512
   sin[421]  =  16'b1101111000011000;     //421pi/512
   cos[421]  =  16'b1100100110111000;     //421pi/512
   sin[422]  =  16'b1101111001101101;     //422pi/512
   cos[422]  =  16'b1100100110000011;     //422pi/512
   sin[423]  =  16'b1101111011000011;     //423pi/512
   cos[423]  =  16'b1100100101001111;     //423pi/512
   sin[424]  =  16'b1101111100011001;     //424pi/512
   cos[424]  =  16'b1100100100011011;     //424pi/512
   sin[425]  =  16'b1101111101101111;     //425pi/512
   cos[425]  =  16'b1100100011101000;     //425pi/512
   sin[426]  =  16'b1101111111000110;     //426pi/512
   cos[426]  =  16'b1100100010110101;     //426pi/512
   sin[427]  =  16'b1110000000011101;     //427pi/512
   cos[427]  =  16'b1100100010000010;     //427pi/512
   sin[428]  =  16'b1110000001110100;     //428pi/512
   cos[428]  =  16'b1100100001010000;     //428pi/512
   sin[429]  =  16'b1110000011001100;     //429pi/512
   cos[429]  =  16'b1100100000011111;     //429pi/512
   sin[430]  =  16'b1110000100100100;     //430pi/512
   cos[430]  =  16'b1100011111101110;     //430pi/512
   sin[431]  =  16'b1110000101111100;     //431pi/512
   cos[431]  =  16'b1100011110111110;     //431pi/512
   sin[432]  =  16'b1110000111010101;     //432pi/512
   cos[432]  =  16'b1100011110001111;     //432pi/512
   sin[433]  =  16'b1110001000101101;     //433pi/512
   cos[433]  =  16'b1100011101011111;     //433pi/512
   sin[434]  =  16'b1110001010000111;     //434pi/512
   cos[434]  =  16'b1100011100110001;     //434pi/512
   sin[435]  =  16'b1110001011100000;     //435pi/512
   cos[435]  =  16'b1100011100000011;     //435pi/512
   sin[436]  =  16'b1110001100111010;     //436pi/512
   cos[436]  =  16'b1100011011010101;     //436pi/512
   sin[437]  =  16'b1110001110010100;     //437pi/512
   cos[437]  =  16'b1100011010101000;     //437pi/512
   sin[438]  =  16'b1110001111101110;     //438pi/512
   cos[438]  =  16'b1100011001111100;     //438pi/512
   sin[439]  =  16'b1110010001001000;     //439pi/512
   cos[439]  =  16'b1100011001010000;     //439pi/512
   sin[440]  =  16'b1110010010100011;     //440pi/512
   cos[440]  =  16'b1100011000100101;     //440pi/512
   sin[441]  =  16'b1110010011111110;     //441pi/512
   cos[441]  =  16'b1100010111111010;     //441pi/512
   sin[442]  =  16'b1110010101011001;     //442pi/512
   cos[442]  =  16'b1100010111010000;     //442pi/512
   sin[443]  =  16'b1110010110110101;     //443pi/512
   cos[443]  =  16'b1100010110100111;     //443pi/512
   sin[444]  =  16'b1110011000010001;     //444pi/512
   cos[444]  =  16'b1100010101111110;     //444pi/512
   sin[445]  =  16'b1110011001101101;     //445pi/512
   cos[445]  =  16'b1100010101010101;     //445pi/512
   sin[446]  =  16'b1110011011001001;     //446pi/512
   cos[446]  =  16'b1100010100101101;     //446pi/512
   sin[447]  =  16'b1110011100100101;     //447pi/512
   cos[447]  =  16'b1100010100000110;     //447pi/512
   sin[448]  =  16'b1110011110000010;     //448pi/512
   cos[448]  =  16'b1100010011011111;     //448pi/512
   sin[449]  =  16'b1110011111011111;     //449pi/512
   cos[449]  =  16'b1100010010111001;     //449pi/512
   sin[450]  =  16'b1110100000111100;     //450pi/512
   cos[450]  =  16'b1100010010010011;     //450pi/512
   sin[451]  =  16'b1110100010011010;     //451pi/512
   cos[451]  =  16'b1100010001101110;     //451pi/512
   sin[452]  =  16'b1110100011110111;     //452pi/512
   cos[452]  =  16'b1100010001001010;     //452pi/512
   sin[453]  =  16'b1110100101010101;     //453pi/512
   cos[453]  =  16'b1100010000100110;     //453pi/512
   sin[454]  =  16'b1110100110110100;     //454pi/512
   cos[454]  =  16'b1100010000000011;     //454pi/512
   sin[455]  =  16'b1110101000010010;     //455pi/512
   cos[455]  =  16'b1100001111100000;     //455pi/512
   sin[456]  =  16'b1110101001110000;     //456pi/512
   cos[456]  =  16'b1100001110111110;     //456pi/512
   sin[457]  =  16'b1110101011001111;     //457pi/512
   cos[457]  =  16'b1100001110011100;     //457pi/512
   sin[458]  =  16'b1110101100101110;     //458pi/512
   cos[458]  =  16'b1100001101111011;     //458pi/512
   sin[459]  =  16'b1110101110001101;     //459pi/512
   cos[459]  =  16'b1100001101011011;     //459pi/512
   sin[460]  =  16'b1110101111101101;     //460pi/512
   cos[460]  =  16'b1100001100111011;     //460pi/512
   sin[461]  =  16'b1110110001001100;     //461pi/512
   cos[461]  =  16'b1100001100011100;     //461pi/512
   sin[462]  =  16'b1110110010101100;     //462pi/512
   cos[462]  =  16'b1100001011111101;     //462pi/512
   sin[463]  =  16'b1110110100001100;     //463pi/512
   cos[463]  =  16'b1100001011011111;     //463pi/512
   sin[464]  =  16'b1110110101101100;     //464pi/512
   cos[464]  =  16'b1100001011000001;     //464pi/512
   sin[465]  =  16'b1110110111001100;     //465pi/512
   cos[465]  =  16'b1100001010100101;     //465pi/512
   sin[466]  =  16'b1110111000101101;     //466pi/512
   cos[466]  =  16'b1100001010001000;     //466pi/512
   sin[467]  =  16'b1110111010001101;     //467pi/512
   cos[467]  =  16'b1100001001101101;     //467pi/512
   sin[468]  =  16'b1110111011101110;     //468pi/512
   cos[468]  =  16'b1100001001010001;     //468pi/512
   sin[469]  =  16'b1110111101001111;     //469pi/512
   cos[469]  =  16'b1100001000110111;     //469pi/512
   sin[470]  =  16'b1110111110110000;     //470pi/512
   cos[470]  =  16'b1100001000011101;     //470pi/512
   sin[471]  =  16'b1111000000010010;     //471pi/512
   cos[471]  =  16'b1100001000000100;     //471pi/512
   sin[472]  =  16'b1111000001110011;     //472pi/512
   cos[472]  =  16'b1100000111101011;     //472pi/512
   sin[473]  =  16'b1111000011010101;     //473pi/512
   cos[473]  =  16'b1100000111010011;     //473pi/512
   sin[474]  =  16'b1111000100110110;     //474pi/512
   cos[474]  =  16'b1100000110111011;     //474pi/512
   sin[475]  =  16'b1111000110011000;     //475pi/512
   cos[475]  =  16'b1100000110100100;     //475pi/512
   sin[476]  =  16'b1111000111111010;     //476pi/512
   cos[476]  =  16'b1100000110001110;     //476pi/512
   sin[477]  =  16'b1111001001011100;     //477pi/512
   cos[477]  =  16'b1100000101111000;     //477pi/512
   sin[478]  =  16'b1111001010111111;     //478pi/512
   cos[478]  =  16'b1100000101100011;     //478pi/512
   sin[479]  =  16'b1111001100100001;     //479pi/512
   cos[479]  =  16'b1100000101001111;     //479pi/512
   sin[480]  =  16'b1111001110000100;     //480pi/512
   cos[480]  =  16'b1100000100111011;     //480pi/512
   sin[481]  =  16'b1111001111100110;     //481pi/512
   cos[481]  =  16'b1100000100101000;     //481pi/512
   sin[482]  =  16'b1111010001001001;     //482pi/512
   cos[482]  =  16'b1100000100010101;     //482pi/512
   sin[483]  =  16'b1111010010101100;     //483pi/512
   cos[483]  =  16'b1100000100000011;     //483pi/512
   sin[484]  =  16'b1111010100001111;     //484pi/512
   cos[484]  =  16'b1100000011110001;     //484pi/512
   sin[485]  =  16'b1111010101110010;     //485pi/512
   cos[485]  =  16'b1100000011100000;     //485pi/512
   sin[486]  =  16'b1111010111010101;     //486pi/512
   cos[486]  =  16'b1100000011010000;     //486pi/512
   sin[487]  =  16'b1111011000111001;     //487pi/512
   cos[487]  =  16'b1100000011000000;     //487pi/512
   sin[488]  =  16'b1111011010011100;     //488pi/512
   cos[488]  =  16'b1100000010110001;     //488pi/512
   sin[489]  =  16'b1111011011111111;     //489pi/512
   cos[489]  =  16'b1100000010100011;     //489pi/512
   sin[490]  =  16'b1111011101100011;     //490pi/512
   cos[490]  =  16'b1100000010010101;     //490pi/512
   sin[491]  =  16'b1111011111000111;     //491pi/512
   cos[491]  =  16'b1100000010001000;     //491pi/512
   sin[492]  =  16'b1111100000101010;     //492pi/512
   cos[492]  =  16'b1100000001111011;     //492pi/512
   sin[493]  =  16'b1111100010001110;     //493pi/512
   cos[493]  =  16'b1100000001101111;     //493pi/512
   sin[494]  =  16'b1111100011110010;     //494pi/512
   cos[494]  =  16'b1100000001100100;     //494pi/512
   sin[495]  =  16'b1111100101010110;     //495pi/512
   cos[495]  =  16'b1100000001011001;     //495pi/512
   sin[496]  =  16'b1111100110111010;     //496pi/512
   cos[496]  =  16'b1100000001001111;     //496pi/512
   sin[497]  =  16'b1111101000011110;     //497pi/512
   cos[497]  =  16'b1100000001000101;     //497pi/512
   sin[498]  =  16'b1111101010000010;     //498pi/512
   cos[498]  =  16'b1100000000111100;     //498pi/512
   sin[499]  =  16'b1111101011100110;     //499pi/512
   cos[499]  =  16'b1100000000110100;     //499pi/512
   sin[500]  =  16'b1111101101001011;     //500pi/512
   cos[500]  =  16'b1100000000101100;     //500pi/512
   sin[501]  =  16'b1111101110101111;     //501pi/512
   cos[501]  =  16'b1100000000100101;     //501pi/512
   sin[502]  =  16'b1111110000010011;     //502pi/512
   cos[502]  =  16'b1100000000011111;     //502pi/512
   sin[503]  =  16'b1111110001111000;     //503pi/512
   cos[503]  =  16'b1100000000011001;     //503pi/512
   sin[504]  =  16'b1111110011011100;     //504pi/512
   cos[504]  =  16'b1100000000010100;     //504pi/512
   sin[505]  =  16'b1111110101000000;     //505pi/512
   cos[505]  =  16'b1100000000001111;     //505pi/512
   sin[506]  =  16'b1111110110100101;     //506pi/512
   cos[506]  =  16'b1100000000001011;     //506pi/512
   sin[507]  =  16'b1111111000001001;     //507pi/512
   cos[507]  =  16'b1100000000001000;     //507pi/512
   sin[508]  =  16'b1111111001101110;     //508pi/512
   cos[508]  =  16'b1100000000000101;     //508pi/512
   sin[509]  =  16'b1111111011010010;     //509pi/512
   cos[509]  =  16'b1100000000000011;     //509pi/512
   sin[510]  =  16'b1111111100110111;     //510pi/512
   cos[510]  =  16'b1100000000000001;     //510pi/512
   sin[511]  =  16'b1111111110011011;     //511pi/512
   cos[511]  =  16'b1100000000000000;     //511pi/512
   m_sin[0]  =  16'b0000000000000000;     //0pi/512
   m_cos[0]  =  16'b0100000000000000;     //0pi/512
   m_sin[1]  =  16'b1111111110100000;     //1pi/512
   m_cos[1]  =  16'b0011111111111111;     //1pi/512
   m_sin[2]  =  16'b1111111101000001;     //2pi/512
   m_cos[2]  =  16'b0011111111111110;     //2pi/512
   m_sin[3]  =  16'b1111111011100010;     //3pi/512
   m_cos[3]  =  16'b0011111111111101;     //3pi/512
   m_sin[4]  =  16'b1111111010000010;     //4pi/512
   m_cos[4]  =  16'b0011111111111011;     //4pi/512
   m_sin[5]  =  16'b1111111000100011;     //5pi/512
   m_cos[5]  =  16'b0011111111111001;     //5pi/512
   m_sin[6]  =  16'b1111110111000011;     //6pi/512
   m_cos[6]  =  16'b0011111111110101;     //6pi/512
   m_sin[7]  =  16'b1111110101100100;     //7pi/512
   m_cos[7]  =  16'b0011111111110010;     //7pi/512
   m_sin[8]  =  16'b1111110100000100;     //8pi/512
   m_cos[8]  =  16'b0011111111101110;     //8pi/512
   m_sin[9]  =  16'b1111110010100101;     //9pi/512
   m_cos[9]  =  16'b0011111111101001;     //9pi/512
   m_sin[10]  =  16'b1111110001000101;     //10pi/512
   m_cos[10]  =  16'b0011111111100100;     //10pi/512
   m_sin[11]  =  16'b1111101111100110;     //11pi/512
   m_cos[11]  =  16'b0011111111011110;     //11pi/512
   m_sin[12]  =  16'b1111101110000111;     //12pi/512
   m_cos[12]  =  16'b0011111111010111;     //12pi/512
   m_sin[13]  =  16'b1111101100101000;     //13pi/512
   m_cos[13]  =  16'b0011111111010000;     //13pi/512
   m_sin[14]  =  16'b1111101011001000;     //14pi/512
   m_cos[14]  =  16'b0011111111001001;     //14pi/512
   m_sin[15]  =  16'b1111101001101001;     //15pi/512
   m_cos[15]  =  16'b0011111111000001;     //15pi/512
   m_sin[16]  =  16'b1111101000001010;     //16pi/512
   m_cos[16]  =  16'b0011111110111000;     //16pi/512
   m_sin[17]  =  16'b1111100110101011;     //17pi/512
   m_cos[17]  =  16'b0011111110101111;     //17pi/512
   m_sin[18]  =  16'b1111100101001100;     //18pi/512
   m_cos[18]  =  16'b0011111110100101;     //18pi/512
   m_sin[19]  =  16'b1111100011101101;     //19pi/512
   m_cos[19]  =  16'b0011111110011011;     //19pi/512
   m_sin[20]  =  16'b1111100010001110;     //20pi/512
   m_cos[20]  =  16'b0011111110010000;     //20pi/512
   m_sin[21]  =  16'b1111100000101111;     //21pi/512
   m_cos[21]  =  16'b0011111110000101;     //21pi/512
   m_sin[22]  =  16'b1111011111010001;     //22pi/512
   m_cos[22]  =  16'b0011111101111001;     //22pi/512
   m_sin[23]  =  16'b1111011101110010;     //23pi/512
   m_cos[23]  =  16'b0011111101101100;     //23pi/512
   m_sin[24]  =  16'b1111011100010011;     //24pi/512
   m_cos[24]  =  16'b0011111101011111;     //24pi/512
   m_sin[25]  =  16'b1111011010110101;     //25pi/512
   m_cos[25]  =  16'b0011111101010010;     //25pi/512
   m_sin[26]  =  16'b1111011001010110;     //26pi/512
   m_cos[26]  =  16'b0011111101000100;     //26pi/512
   m_sin[27]  =  16'b1111010111111000;     //27pi/512
   m_cos[27]  =  16'b0011111100110101;     //27pi/512
   m_sin[28]  =  16'b1111010110011010;     //28pi/512
   m_cos[28]  =  16'b0011111100100110;     //28pi/512
   m_sin[29]  =  16'b1111010100111100;     //29pi/512
   m_cos[29]  =  16'b0011111100010110;     //29pi/512
   m_sin[30]  =  16'b1111010011011101;     //30pi/512
   m_cos[30]  =  16'b0011111100000110;     //30pi/512
   m_sin[31]  =  16'b1111010001111111;     //31pi/512
   m_cos[31]  =  16'b0011111011110101;     //31pi/512
   m_sin[32]  =  16'b1111010000100010;     //32pi/512
   m_cos[32]  =  16'b0011111011100011;     //32pi/512
   m_sin[33]  =  16'b1111001111000100;     //33pi/512
   m_cos[33]  =  16'b0011111011010001;     //33pi/512
   m_sin[34]  =  16'b1111001101100110;     //34pi/512
   m_cos[34]  =  16'b0011111010111111;     //34pi/512
   m_sin[35]  =  16'b1111001100001000;     //35pi/512
   m_cos[35]  =  16'b0011111010101100;     //35pi/512
   m_sin[36]  =  16'b1111001010101011;     //36pi/512
   m_cos[36]  =  16'b0011111010011000;     //36pi/512
   m_sin[37]  =  16'b1111001001001110;     //37pi/512
   m_cos[37]  =  16'b0011111010000100;     //37pi/512
   m_sin[38]  =  16'b1111000111110000;     //38pi/512
   m_cos[38]  =  16'b0011111001101111;     //38pi/512
   m_sin[39]  =  16'b1111000110010011;     //39pi/512
   m_cos[39]  =  16'b0011111001011010;     //39pi/512
   m_sin[40]  =  16'b1111000100110110;     //40pi/512
   m_cos[40]  =  16'b0011111001000100;     //40pi/512
   m_sin[41]  =  16'b1111000011011001;     //41pi/512
   m_cos[41]  =  16'b0011111000101110;     //41pi/512
   m_sin[42]  =  16'b1111000001111101;     //42pi/512
   m_cos[42]  =  16'b0011111000010111;     //42pi/512
   m_sin[43]  =  16'b1111000000100000;     //43pi/512
   m_cos[43]  =  16'b0011111000000000;     //43pi/512
   m_sin[44]  =  16'b1110111111000100;     //44pi/512
   m_cos[44]  =  16'b0011110111101000;     //44pi/512
   m_sin[45]  =  16'b1110111101100111;     //45pi/512
   m_cos[45]  =  16'b0011110111001111;     //45pi/512
   m_sin[46]  =  16'b1110111100001011;     //46pi/512
   m_cos[46]  =  16'b0011110110110110;     //46pi/512
   m_sin[47]  =  16'b1110111010101111;     //47pi/512
   m_cos[47]  =  16'b0011110110011100;     //47pi/512
   m_sin[48]  =  16'b1110111001010011;     //48pi/512
   m_cos[48]  =  16'b0011110110000010;     //48pi/512
   m_sin[49]  =  16'b1110110111111000;     //49pi/512
   m_cos[49]  =  16'b0011110101101000;     //49pi/512
   m_sin[50]  =  16'b1110110110011100;     //50pi/512
   m_cos[50]  =  16'b0011110101001101;     //50pi/512
   m_sin[51]  =  16'b1110110101000001;     //51pi/512
   m_cos[51]  =  16'b0011110100110001;     //51pi/512
   m_sin[52]  =  16'b1110110011100101;     //52pi/512
   m_cos[52]  =  16'b0011110100010101;     //52pi/512
   m_sin[53]  =  16'b1110110010001010;     //53pi/512
   m_cos[53]  =  16'b0011110011111000;     //53pi/512
   m_sin[54]  =  16'b1110110000110000;     //54pi/512
   m_cos[54]  =  16'b0011110011011011;     //54pi/512
   m_sin[55]  =  16'b1110101111010101;     //55pi/512
   m_cos[55]  =  16'b0011110010111101;     //55pi/512
   m_sin[56]  =  16'b1110101101111010;     //56pi/512
   m_cos[56]  =  16'b0011110010011110;     //56pi/512
   m_sin[57]  =  16'b1110101100100000;     //57pi/512
   m_cos[57]  =  16'b0011110001111111;     //57pi/512
   m_sin[58]  =  16'b1110101011000110;     //58pi/512
   m_cos[58]  =  16'b0011110001100000;     //58pi/512
   m_sin[59]  =  16'b1110101001101100;     //59pi/512
   m_cos[59]  =  16'b0011110001000000;     //59pi/512
   m_sin[60]  =  16'b1110101000010010;     //60pi/512
   m_cos[60]  =  16'b0011110000100000;     //60pi/512
   m_sin[61]  =  16'b1110100110111000;     //61pi/512
   m_cos[61]  =  16'b0011101111111111;     //61pi/512
   m_sin[62]  =  16'b1110100101011111;     //62pi/512
   m_cos[62]  =  16'b0011101111011101;     //62pi/512
   m_sin[63]  =  16'b1110100100000110;     //63pi/512
   m_cos[63]  =  16'b0011101110111011;     //63pi/512
   m_sin[64]  =  16'b1110100010101101;     //64pi/512
   m_cos[64]  =  16'b0011101110011001;     //64pi/512
   m_sin[65]  =  16'b1110100001010100;     //65pi/512
   m_cos[65]  =  16'b0011101101110101;     //65pi/512
   m_sin[66]  =  16'b1110011111111011;     //66pi/512
   m_cos[66]  =  16'b0011101101010010;     //66pi/512
   m_sin[67]  =  16'b1110011110100011;     //67pi/512
   m_cos[67]  =  16'b0011101100101110;     //67pi/512
   m_sin[68]  =  16'b1110011101001010;     //68pi/512
   m_cos[68]  =  16'b0011101100001001;     //68pi/512
   m_sin[69]  =  16'b1110011011110010;     //69pi/512
   m_cos[69]  =  16'b0011101011100100;     //69pi/512
   m_sin[70]  =  16'b1110011010011011;     //70pi/512
   m_cos[70]  =  16'b0011101010111110;     //70pi/512
   m_sin[71]  =  16'b1110011001000011;     //71pi/512
   m_cos[71]  =  16'b0011101010011000;     //71pi/512
   m_sin[72]  =  16'b1110010111101100;     //72pi/512
   m_cos[72]  =  16'b0011101001110010;     //72pi/512
   m_sin[73]  =  16'b1110010110010101;     //73pi/512
   m_cos[73]  =  16'b0011101001001010;     //73pi/512
   m_sin[74]  =  16'b1110010100111110;     //74pi/512
   m_cos[74]  =  16'b0011101000100011;     //74pi/512
   m_sin[75]  =  16'b1110010011100111;     //75pi/512
   m_cos[75]  =  16'b0011100111111011;     //75pi/512
   m_sin[76]  =  16'b1110010010010001;     //76pi/512
   m_cos[76]  =  16'b0011100111010010;     //76pi/512
   m_sin[77]  =  16'b1110010000111011;     //77pi/512
   m_cos[77]  =  16'b0011100110101001;     //77pi/512
   m_sin[78]  =  16'b1110001111100101;     //78pi/512
   m_cos[78]  =  16'b0011100101111111;     //78pi/512
   m_sin[79]  =  16'b1110001110001111;     //79pi/512
   m_cos[79]  =  16'b0011100101010101;     //79pi/512
   m_sin[80]  =  16'b1110001100111010;     //80pi/512
   m_cos[80]  =  16'b0011100100101010;     //80pi/512
   m_sin[81]  =  16'b1110001011100100;     //81pi/512
   m_cos[81]  =  16'b0011100011111111;     //81pi/512
   m_sin[82]  =  16'b1110001010001111;     //82pi/512
   m_cos[82]  =  16'b0011100011010011;     //82pi/512
   m_sin[83]  =  16'b1110001000111011;     //83pi/512
   m_cos[83]  =  16'b0011100010100111;     //83pi/512
   m_sin[84]  =  16'b1110000111100110;     //84pi/512
   m_cos[84]  =  16'b0011100001111010;     //84pi/512
   m_sin[85]  =  16'b1110000110010010;     //85pi/512
   m_cos[85]  =  16'b0011100001001101;     //85pi/512
   m_sin[86]  =  16'b1110000100111110;     //86pi/512
   m_cos[86]  =  16'b0011100000100000;     //86pi/512
   m_sin[87]  =  16'b1110000011101011;     //87pi/512
   m_cos[87]  =  16'b0011011111110001;     //87pi/512
   m_sin[88]  =  16'b1110000010010111;     //88pi/512
   m_cos[88]  =  16'b0011011111000011;     //88pi/512
   m_sin[89]  =  16'b1110000001000100;     //89pi/512
   m_cos[89]  =  16'b0011011110010100;     //89pi/512
   m_sin[90]  =  16'b1101111111110001;     //90pi/512
   m_cos[90]  =  16'b0011011101100100;     //90pi/512
   m_sin[91]  =  16'b1101111110011111;     //91pi/512
   m_cos[91]  =  16'b0011011100110100;     //91pi/512
   m_sin[92]  =  16'b1101111101001101;     //92pi/512
   m_cos[92]  =  16'b0011011100000011;     //92pi/512
   m_sin[93]  =  16'b1101111011111011;     //93pi/512
   m_cos[93]  =  16'b0011011011010010;     //93pi/512
   m_sin[94]  =  16'b1101111010101001;     //94pi/512
   m_cos[94]  =  16'b0011011010100001;     //94pi/512
   m_sin[95]  =  16'b1101111001011000;     //95pi/512
   m_cos[95]  =  16'b0011011001101111;     //95pi/512
   m_sin[96]  =  16'b1101111000000111;     //96pi/512
   m_cos[96]  =  16'b0011011000111100;     //96pi/512
   m_sin[97]  =  16'b1101110110110110;     //97pi/512
   m_cos[97]  =  16'b0011011000001010;     //97pi/512
   m_sin[98]  =  16'b1101110101100101;     //98pi/512
   m_cos[98]  =  16'b0011010111010110;     //98pi/512
   m_sin[99]  =  16'b1101110100010101;     //99pi/512
   m_cos[99]  =  16'b0011010110100010;     //99pi/512
   m_sin[100]  =  16'b1101110011000101;     //100pi/512
   m_cos[100]  =  16'b0011010101101110;     //100pi/512
   m_sin[101]  =  16'b1101110001110110;     //101pi/512
   m_cos[101]  =  16'b0011010100111001;     //101pi/512
   m_sin[102]  =  16'b1101110000100110;     //102pi/512
   m_cos[102]  =  16'b0011010100000100;     //102pi/512
   m_sin[103]  =  16'b1101101111010111;     //103pi/512
   m_cos[103]  =  16'b0011010011001110;     //103pi/512
   m_sin[104]  =  16'b1101101110001001;     //104pi/512
   m_cos[104]  =  16'b0011010010011000;     //104pi/512
   m_sin[105]  =  16'b1101101100111011;     //105pi/512
   m_cos[105]  =  16'b0011010001100001;     //105pi/512
   m_sin[106]  =  16'b1101101011101101;     //106pi/512
   m_cos[106]  =  16'b0011010000101010;     //106pi/512
   m_sin[107]  =  16'b1101101010011111;     //107pi/512
   m_cos[107]  =  16'b0011001111110011;     //107pi/512
   m_sin[108]  =  16'b1101101001010001;     //108pi/512
   m_cos[108]  =  16'b0011001110111011;     //108pi/512
   m_sin[109]  =  16'b1101101000000100;     //109pi/512
   m_cos[109]  =  16'b0011001110000010;     //109pi/512
   m_sin[110]  =  16'b1101100110111000;     //110pi/512
   m_cos[110]  =  16'b0011001101001001;     //110pi/512
   m_sin[111]  =  16'b1101100101101011;     //111pi/512
   m_cos[111]  =  16'b0011001100010000;     //111pi/512
   m_sin[112]  =  16'b1101100100011111;     //112pi/512
   m_cos[112]  =  16'b0011001011010110;     //112pi/512
   m_sin[113]  =  16'b1101100011010100;     //113pi/512
   m_cos[113]  =  16'b0011001010011100;     //113pi/512
   m_sin[114]  =  16'b1101100010001000;     //114pi/512
   m_cos[114]  =  16'b0011001001100001;     //114pi/512
   m_sin[115]  =  16'b1101100000111101;     //115pi/512
   m_cos[115]  =  16'b0011001000100110;     //115pi/512
   m_sin[116]  =  16'b1101011111110011;     //116pi/512
   m_cos[116]  =  16'b0011000111101011;     //116pi/512
   m_sin[117]  =  16'b1101011110101000;     //117pi/512
   m_cos[117]  =  16'b0011000110101111;     //117pi/512
   m_sin[118]  =  16'b1101011101011110;     //118pi/512
   m_cos[118]  =  16'b0011000101110010;     //118pi/512
   m_sin[119]  =  16'b1101011100010101;     //119pi/512
   m_cos[119]  =  16'b0011000100110101;     //119pi/512
   m_sin[120]  =  16'b1101011011001011;     //120pi/512
   m_cos[120]  =  16'b0011000011111000;     //120pi/512
   m_sin[121]  =  16'b1101011010000011;     //121pi/512
   m_cos[121]  =  16'b0011000010111010;     //121pi/512
   m_sin[122]  =  16'b1101011000111010;     //122pi/512
   m_cos[122]  =  16'b0011000001111100;     //122pi/512
   m_sin[123]  =  16'b1101010111110010;     //123pi/512
   m_cos[123]  =  16'b0011000000111110;     //123pi/512
   m_sin[124]  =  16'b1101010110101010;     //124pi/512
   m_cos[124]  =  16'b0010111111111111;     //124pi/512
   m_sin[125]  =  16'b1101010101100011;     //125pi/512
   m_cos[125]  =  16'b0010111110111111;     //125pi/512
   m_sin[126]  =  16'b1101010100011100;     //126pi/512
   m_cos[126]  =  16'b0010111101111111;     //126pi/512
   m_sin[127]  =  16'b1101010011010101;     //127pi/512
   m_cos[127]  =  16'b0010111100111111;     //127pi/512
   m_sin[128]  =  16'b1101010010001111;     //128pi/512
   m_cos[128]  =  16'b0010111011111111;     //128pi/512
   m_sin[129]  =  16'b1101010001001001;     //129pi/512
   m_cos[129]  =  16'b0010111010111110;     //129pi/512
   m_sin[130]  =  16'b1101010000000011;     //130pi/512
   m_cos[130]  =  16'b0010111001111100;     //130pi/512
   m_sin[131]  =  16'b1101001110111110;     //131pi/512
   m_cos[131]  =  16'b0010111000111010;     //131pi/512
   m_sin[132]  =  16'b1101001101111001;     //132pi/512
   m_cos[132]  =  16'b0010110111111000;     //132pi/512
   m_sin[133]  =  16'b1101001100110101;     //133pi/512
   m_cos[133]  =  16'b0010110110110101;     //133pi/512
   m_sin[134]  =  16'b1101001011110001;     //134pi/512
   m_cos[134]  =  16'b0010110101110010;     //134pi/512
   m_sin[135]  =  16'b1101001010101101;     //135pi/512
   m_cos[135]  =  16'b0010110100101111;     //135pi/512
   m_sin[136]  =  16'b1101001001101010;     //136pi/512
   m_cos[136]  =  16'b0010110011101011;     //136pi/512
   m_sin[137]  =  16'b1101001000100111;     //137pi/512
   m_cos[137]  =  16'b0010110010100111;     //137pi/512
   m_sin[138]  =  16'b1101000111100101;     //138pi/512
   m_cos[138]  =  16'b0010110001100010;     //138pi/512
   m_sin[139]  =  16'b1101000110100010;     //139pi/512
   m_cos[139]  =  16'b0010110000011101;     //139pi/512
   m_sin[140]  =  16'b1101000101100001;     //140pi/512
   m_cos[140]  =  16'b0010101111011000;     //140pi/512
   m_sin[141]  =  16'b1101000100100000;     //141pi/512
   m_cos[141]  =  16'b0010101110010010;     //141pi/512
   m_sin[142]  =  16'b1101000011011111;     //142pi/512
   m_cos[142]  =  16'b0010101101001100;     //142pi/512
   m_sin[143]  =  16'b1101000010011110;     //143pi/512
   m_cos[143]  =  16'b0010101100000101;     //143pi/512
   m_sin[144]  =  16'b1101000001011110;     //144pi/512
   m_cos[144]  =  16'b0010101010111111;     //144pi/512
   m_sin[145]  =  16'b1101000000011111;     //145pi/512
   m_cos[145]  =  16'b0010101001110111;     //145pi/512
   m_sin[146]  =  16'b1100111111100000;     //146pi/512
   m_cos[146]  =  16'b0010101000110000;     //146pi/512
   m_sin[147]  =  16'b1100111110100001;     //147pi/512
   m_cos[147]  =  16'b0010100111101000;     //147pi/512
   m_sin[148]  =  16'b1100111101100011;     //148pi/512
   m_cos[148]  =  16'b0010100110011111;     //148pi/512
   m_sin[149]  =  16'b1100111100100101;     //149pi/512
   m_cos[149]  =  16'b0010100101010111;     //149pi/512
   m_sin[150]  =  16'b1100111011100111;     //150pi/512
   m_cos[150]  =  16'b0010100100001110;     //150pi/512
   m_sin[151]  =  16'b1100111010101010;     //151pi/512
   m_cos[151]  =  16'b0010100011000100;     //151pi/512
   m_sin[152]  =  16'b1100111001101110;     //152pi/512
   m_cos[152]  =  16'b0010100001111010;     //152pi/512
   m_sin[153]  =  16'b1100111000110001;     //153pi/512
   m_cos[153]  =  16'b0010100000110000;     //153pi/512
   m_sin[154]  =  16'b1100110111110110;     //154pi/512
   m_cos[154]  =  16'b0010011111100110;     //154pi/512
   m_sin[155]  =  16'b1100110110111010;     //155pi/512
   m_cos[155]  =  16'b0010011110011011;     //155pi/512
   m_sin[156]  =  16'b1100110101111111;     //156pi/512
   m_cos[156]  =  16'b0010011101010000;     //156pi/512
   m_sin[157]  =  16'b1100110101000101;     //157pi/512
   m_cos[157]  =  16'b0010011100000100;     //157pi/512
   m_sin[158]  =  16'b1100110100001011;     //158pi/512
   m_cos[158]  =  16'b0010011010111000;     //158pi/512
   m_sin[159]  =  16'b1100110011010001;     //159pi/512
   m_cos[159]  =  16'b0010011001101100;     //159pi/512
   m_sin[160]  =  16'b1100110010011000;     //160pi/512
   m_cos[160]  =  16'b0010011000011111;     //160pi/512
   m_sin[161]  =  16'b1100110001100000;     //161pi/512
   m_cos[161]  =  16'b0010010111010011;     //161pi/512
   m_sin[162]  =  16'b1100110000100111;     //162pi/512
   m_cos[162]  =  16'b0010010110000101;     //162pi/512
   m_sin[163]  =  16'b1100101111110000;     //163pi/512
   m_cos[163]  =  16'b0010010100111000;     //163pi/512
   m_sin[164]  =  16'b1100101110111000;     //164pi/512
   m_cos[164]  =  16'b0010010011101010;     //164pi/512
   m_sin[165]  =  16'b1100101110000001;     //165pi/512
   m_cos[165]  =  16'b0010010010011100;     //165pi/512
   m_sin[166]  =  16'b1100101101001011;     //166pi/512
   m_cos[166]  =  16'b0010010001001101;     //166pi/512
   m_sin[167]  =  16'b1100101100010101;     //167pi/512
   m_cos[167]  =  16'b0010001111111110;     //167pi/512
   m_sin[168]  =  16'b1100101011100000;     //168pi/512
   m_cos[168]  =  16'b0010001110101111;     //168pi/512
   m_sin[169]  =  16'b1100101010101011;     //169pi/512
   m_cos[169]  =  16'b0010001101100000;     //169pi/512
   m_sin[170]  =  16'b1100101001110110;     //170pi/512
   m_cos[170]  =  16'b0010001100010000;     //170pi/512
   m_sin[171]  =  16'b1100101001000010;     //171pi/512
   m_cos[171]  =  16'b0010001011000000;     //171pi/512
   m_sin[172]  =  16'b1100101000001110;     //172pi/512
   m_cos[172]  =  16'b0010001001110000;     //172pi/512
   m_sin[173]  =  16'b1100100111011011;     //173pi/512
   m_cos[173]  =  16'b0010001000011111;     //173pi/512
   m_sin[174]  =  16'b1100100110101000;     //174pi/512
   m_cos[174]  =  16'b0010000111001110;     //174pi/512
   m_sin[175]  =  16'b1100100101110110;     //175pi/512
   m_cos[175]  =  16'b0010000101111101;     //175pi/512
   m_sin[176]  =  16'b1100100101000100;     //176pi/512
   m_cos[176]  =  16'b0010000100101011;     //176pi/512
   m_sin[177]  =  16'b1100100100010011;     //177pi/512
   m_cos[177]  =  16'b0010000011011010;     //177pi/512
   m_sin[178]  =  16'b1100100011100010;     //178pi/512
   m_cos[178]  =  16'b0010000010001000;     //178pi/512
   m_sin[179]  =  16'b1100100010110010;     //179pi/512
   m_cos[179]  =  16'b0010000000110101;     //179pi/512
   m_sin[180]  =  16'b1100100010000010;     //180pi/512
   m_cos[180]  =  16'b0001111111100010;     //180pi/512
   m_sin[181]  =  16'b1100100001010011;     //181pi/512
   m_cos[181]  =  16'b0001111110010000;     //181pi/512
   m_sin[182]  =  16'b1100100000100100;     //182pi/512
   m_cos[182]  =  16'b0001111100111100;     //182pi/512
   m_sin[183]  =  16'b1100011111110110;     //183pi/512
   m_cos[183]  =  16'b0001111011101001;     //183pi/512
   m_sin[184]  =  16'b1100011111001000;     //184pi/512
   m_cos[184]  =  16'b0001111010010101;     //184pi/512
   m_sin[185]  =  16'b1100011110011010;     //185pi/512
   m_cos[185]  =  16'b0001111001000001;     //185pi/512
   m_sin[186]  =  16'b1100011101101110;     //186pi/512
   m_cos[186]  =  16'b0001110111101101;     //186pi/512
   m_sin[187]  =  16'b1100011101000001;     //187pi/512
   m_cos[187]  =  16'b0001110110011000;     //187pi/512
   m_sin[188]  =  16'b1100011100010101;     //188pi/512
   m_cos[188]  =  16'b0001110101000011;     //188pi/512
   m_sin[189]  =  16'b1100011011101010;     //189pi/512
   m_cos[189]  =  16'b0001110011101110;     //189pi/512
   m_sin[190]  =  16'b1100011010111111;     //190pi/512
   m_cos[190]  =  16'b0001110010011001;     //190pi/512
   m_sin[191]  =  16'b1100011010010100;     //191pi/512
   m_cos[191]  =  16'b0001110001000011;     //191pi/512
   m_sin[192]  =  16'b1100011001101011;     //192pi/512
   m_cos[192]  =  16'b0001101111101110;     //192pi/512
   m_sin[193]  =  16'b1100011001000001;     //193pi/512
   m_cos[193]  =  16'b0001101110011000;     //193pi/512
   m_sin[194]  =  16'b1100011000011000;     //194pi/512
   m_cos[194]  =  16'b0001101101000001;     //194pi/512
   m_sin[195]  =  16'b1100010111110000;     //195pi/512
   m_cos[195]  =  16'b0001101011101011;     //195pi/512
   m_sin[196]  =  16'b1100010111001000;     //196pi/512
   m_cos[196]  =  16'b0001101010010100;     //196pi/512
   m_sin[197]  =  16'b1100010110100000;     //197pi/512
   m_cos[197]  =  16'b0001101000111101;     //197pi/512
   m_sin[198]  =  16'b1100010101111010;     //198pi/512
   m_cos[198]  =  16'b0001100111100110;     //198pi/512
   m_sin[199]  =  16'b1100010101010011;     //199pi/512
   m_cos[199]  =  16'b0001100110001110;     //199pi/512
   m_sin[200]  =  16'b1100010100101101;     //200pi/512
   m_cos[200]  =  16'b0001100100110111;     //200pi/512
   m_sin[201]  =  16'b1100010100001000;     //201pi/512
   m_cos[201]  =  16'b0001100011011111;     //201pi/512
   m_sin[202]  =  16'b1100010011100011;     //202pi/512
   m_cos[202]  =  16'b0001100010000111;     //202pi/512
   m_sin[203]  =  16'b1100010010111111;     //203pi/512
   m_cos[203]  =  16'b0001100000101110;     //203pi/512
   m_sin[204]  =  16'b1100010010011011;     //204pi/512
   m_cos[204]  =  16'b0001011111010110;     //204pi/512
   m_sin[205]  =  16'b1100010001111000;     //205pi/512
   m_cos[205]  =  16'b0001011101111101;     //205pi/512
   m_sin[206]  =  16'b1100010001010101;     //206pi/512
   m_cos[206]  =  16'b0001011100100100;     //206pi/512
   m_sin[207]  =  16'b1100010000110010;     //207pi/512
   m_cos[207]  =  16'b0001011011001011;     //207pi/512
   m_sin[208]  =  16'b1100010000010001;     //208pi/512
   m_cos[208]  =  16'b0001011001110010;     //208pi/512
   m_sin[209]  =  16'b1100001111101111;     //209pi/512
   m_cos[209]  =  16'b0001011000011000;     //209pi/512
   m_sin[210]  =  16'b1100001111001111;     //210pi/512
   m_cos[210]  =  16'b0001010110111110;     //210pi/512
   m_sin[211]  =  16'b1100001110101111;     //211pi/512
   m_cos[211]  =  16'b0001010101100100;     //211pi/512
   m_sin[212]  =  16'b1100001110001111;     //212pi/512
   m_cos[212]  =  16'b0001010100001010;     //212pi/512
   m_sin[213]  =  16'b1100001101110000;     //213pi/512
   m_cos[213]  =  16'b0001010010110000;     //213pi/512
   m_sin[214]  =  16'b1100001101010001;     //214pi/512
   m_cos[214]  =  16'b0001010001010110;     //214pi/512
   m_sin[215]  =  16'b1100001100110011;     //215pi/512
   m_cos[215]  =  16'b0001001111111011;     //215pi/512
   m_sin[216]  =  16'b1100001100010110;     //216pi/512
   m_cos[216]  =  16'b0001001110100000;     //216pi/512
   m_sin[217]  =  16'b1100001011111000;     //217pi/512
   m_cos[217]  =  16'b0001001101000101;     //217pi/512
   m_sin[218]  =  16'b1100001011011100;     //218pi/512
   m_cos[218]  =  16'b0001001011101010;     //218pi/512
   m_sin[219]  =  16'b1100001011000000;     //219pi/512
   m_cos[219]  =  16'b0001001010001111;     //219pi/512
   m_sin[220]  =  16'b1100001010100101;     //220pi/512
   m_cos[220]  =  16'b0001001000110011;     //220pi/512
   m_sin[221]  =  16'b1100001010001010;     //221pi/512
   m_cos[221]  =  16'b0001000111011000;     //221pi/512
   m_sin[222]  =  16'b1100001001101111;     //222pi/512
   m_cos[222]  =  16'b0001000101111100;     //222pi/512
   m_sin[223]  =  16'b1100001001010110;     //223pi/512
   m_cos[223]  =  16'b0001000100100000;     //223pi/512
   m_sin[224]  =  16'b1100001000111100;     //224pi/512
   m_cos[224]  =  16'b0001000011000100;     //224pi/512
   m_sin[225]  =  16'b1100001000100011;     //225pi/512
   m_cos[225]  =  16'b0001000001101000;     //225pi/512
   m_sin[226]  =  16'b1100001000001011;     //226pi/512
   m_cos[226]  =  16'b0001000000001011;     //226pi/512
   m_sin[227]  =  16'b1100000111110100;     //227pi/512
   m_cos[227]  =  16'b0000111110101111;     //227pi/512
   m_sin[228]  =  16'b1100000111011100;     //228pi/512
   m_cos[228]  =  16'b0000111101010010;     //228pi/512
   m_sin[229]  =  16'b1100000111000110;     //229pi/512
   m_cos[229]  =  16'b0000111011110101;     //229pi/512
   m_sin[230]  =  16'b1100000110110000;     //230pi/512
   m_cos[230]  =  16'b0000111010011000;     //230pi/512
   m_sin[231]  =  16'b1100000110011010;     //231pi/512
   m_cos[231]  =  16'b0000111000111011;     //231pi/512
   m_sin[232]  =  16'b1100000110000101;     //232pi/512
   m_cos[232]  =  16'b0000110111011110;     //232pi/512
   m_sin[233]  =  16'b1100000101110001;     //233pi/512
   m_cos[233]  =  16'b0000110110000001;     //233pi/512
   m_sin[234]  =  16'b1100000101011101;     //234pi/512
   m_cos[234]  =  16'b0000110100100011;     //234pi/512
   m_sin[235]  =  16'b1100000101001010;     //235pi/512
   m_cos[235]  =  16'b0000110011000110;     //235pi/512
   m_sin[236]  =  16'b1100000100110111;     //236pi/512
   m_cos[236]  =  16'b0000110001101000;     //236pi/512
   m_sin[237]  =  16'b1100000100100101;     //237pi/512
   m_cos[237]  =  16'b0000110000001010;     //237pi/512
   m_sin[238]  =  16'b1100000100010011;     //238pi/512
   m_cos[238]  =  16'b0000101110101101;     //238pi/512
   m_sin[239]  =  16'b1100000100000010;     //239pi/512
   m_cos[239]  =  16'b0000101101001111;     //239pi/512
   m_sin[240]  =  16'b1100000011110001;     //240pi/512
   m_cos[240]  =  16'b0000101011110001;     //240pi/512
   m_sin[241]  =  16'b1100000011100001;     //241pi/512
   m_cos[241]  =  16'b0000101010010010;     //241pi/512
   m_sin[242]  =  16'b1100000011010010;     //242pi/512
   m_cos[242]  =  16'b0000101000110100;     //242pi/512
   m_sin[243]  =  16'b1100000011000011;     //243pi/512
   m_cos[243]  =  16'b0000100111010110;     //243pi/512
   m_sin[244]  =  16'b1100000010110100;     //244pi/512
   m_cos[244]  =  16'b0000100101110111;     //244pi/512
   m_sin[245]  =  16'b1100000010100110;     //245pi/512
   m_cos[245]  =  16'b0000100100011001;     //245pi/512
   m_sin[246]  =  16'b1100000010011001;     //246pi/512
   m_cos[246]  =  16'b0000100010111010;     //246pi/512
   m_sin[247]  =  16'b1100000010001100;     //247pi/512
   m_cos[247]  =  16'b0000100001011100;     //247pi/512
   m_sin[248]  =  16'b1100000010000000;     //248pi/512
   m_cos[248]  =  16'b0000011111111101;     //248pi/512
   m_sin[249]  =  16'b1100000001110101;     //249pi/512
   m_cos[249]  =  16'b0000011110011110;     //249pi/512
   m_sin[250]  =  16'b1100000001101001;     //250pi/512
   m_cos[250]  =  16'b0000011100111111;     //250pi/512
   m_sin[251]  =  16'b1100000001011111;     //251pi/512
   m_cos[251]  =  16'b0000011011100000;     //251pi/512
   m_sin[252]  =  16'b1100000001010101;     //252pi/512
   m_cos[252]  =  16'b0000011010000001;     //252pi/512
   m_sin[253]  =  16'b1100000001001011;     //253pi/512
   m_cos[253]  =  16'b0000011000100010;     //253pi/512
   m_sin[254]  =  16'b1100000001000011;     //254pi/512
   m_cos[254]  =  16'b0000010111000011;     //254pi/512
   m_sin[255]  =  16'b1100000000111010;     //255pi/512
   m_cos[255]  =  16'b0000010101100100;     //255pi/512
   m_sin[256]  =  16'b1100000000110011;     //256pi/512
   m_cos[256]  =  16'b0000010100000101;     //256pi/512
   m_sin[257]  =  16'b1100000000101011;     //257pi/512
   m_cos[257]  =  16'b0000010010100110;     //257pi/512
   m_sin[258]  =  16'b1100000000100101;     //258pi/512
   m_cos[258]  =  16'b0000010001000110;     //258pi/512
   m_sin[259]  =  16'b1100000000011111;     //259pi/512
   m_cos[259]  =  16'b0000001111100111;     //259pi/512
   m_sin[260]  =  16'b1100000000011001;     //260pi/512
   m_cos[260]  =  16'b0000001110001000;     //260pi/512
   m_sin[261]  =  16'b1100000000010100;     //261pi/512
   m_cos[261]  =  16'b0000001100101000;     //261pi/512
   m_sin[262]  =  16'b1100000000010000;     //262pi/512
   m_cos[262]  =  16'b0000001011001001;     //262pi/512
   m_sin[263]  =  16'b1100000000001100;     //263pi/512
   m_cos[263]  =  16'b0000001001101010;     //263pi/512
   m_sin[264]  =  16'b1100000000001000;     //264pi/512
   m_cos[264]  =  16'b0000001000001010;     //264pi/512
   m_sin[265]  =  16'b1100000000000110;     //265pi/512
   m_cos[265]  =  16'b0000000110101011;     //265pi/512
   m_sin[266]  =  16'b1100000000000011;     //266pi/512
   m_cos[266]  =  16'b0000000101001011;     //266pi/512
   m_sin[267]  =  16'b1100000000000010;     //267pi/512
   m_cos[267]  =  16'b0000000011101100;     //267pi/512
   m_sin[268]  =  16'b1100000000000001;     //268pi/512
   m_cos[268]  =  16'b0000000010001100;     //268pi/512
   m_sin[269]  =  16'b1100000000000000;     //269pi/512
   m_cos[269]  =  16'b0000000000101101;     //269pi/512
   m_sin[270]  =  16'b1100000000000000;     //270pi/512
   m_cos[270]  =  16'b1111111111001110;     //270pi/512
   m_sin[271]  =  16'b1100000000000001;     //271pi/512
   m_cos[271]  =  16'b1111111101101110;     //271pi/512
   m_sin[272]  =  16'b1100000000000010;     //272pi/512
   m_cos[272]  =  16'b1111111100001111;     //272pi/512
   m_sin[273]  =  16'b1100000000000011;     //273pi/512
   m_cos[273]  =  16'b1111111010101111;     //273pi/512
   m_sin[274]  =  16'b1100000000000110;     //274pi/512
   m_cos[274]  =  16'b1111111001010000;     //274pi/512
   m_sin[275]  =  16'b1100000000001001;     //275pi/512
   m_cos[275]  =  16'b1111110111110000;     //275pi/512
   m_sin[276]  =  16'b1100000000001100;     //276pi/512
   m_cos[276]  =  16'b1111110110010001;     //276pi/512
   m_sin[277]  =  16'b1100000000010000;     //277pi/512
   m_cos[277]  =  16'b1111110100110001;     //277pi/512
   m_sin[278]  =  16'b1100000000010100;     //278pi/512
   m_cos[278]  =  16'b1111110011010010;     //278pi/512
   m_sin[279]  =  16'b1100000000011001;     //279pi/512
   m_cos[279]  =  16'b1111110001110011;     //279pi/512
   m_sin[280]  =  16'b1100000000011111;     //280pi/512
   m_cos[280]  =  16'b1111110000010011;     //280pi/512
   m_sin[281]  =  16'b1100000000100101;     //281pi/512
   m_cos[281]  =  16'b1111101110110100;     //281pi/512
   m_sin[282]  =  16'b1100000000101100;     //282pi/512
   m_cos[282]  =  16'b1111101101010101;     //282pi/512
   m_sin[283]  =  16'b1100000000110011;     //283pi/512
   m_cos[283]  =  16'b1111101011110110;     //283pi/512
   m_sin[284]  =  16'b1100000000111011;     //284pi/512
   m_cos[284]  =  16'b1111101010010110;     //284pi/512
   m_sin[285]  =  16'b1100000001000011;     //285pi/512
   m_cos[285]  =  16'b1111101000110111;     //285pi/512
   m_sin[286]  =  16'b1100000001001100;     //286pi/512
   m_cos[286]  =  16'b1111100111011000;     //286pi/512
   m_sin[287]  =  16'b1100000001010101;     //287pi/512
   m_cos[287]  =  16'b1111100101111001;     //287pi/512
   m_sin[288]  =  16'b1100000001011111;     //288pi/512
   m_cos[288]  =  16'b1111100100011010;     //288pi/512
   m_sin[289]  =  16'b1100000001101010;     //289pi/512
   m_cos[289]  =  16'b1111100010111011;     //289pi/512
   m_sin[290]  =  16'b1100000001110101;     //290pi/512
   m_cos[290]  =  16'b1111100001011100;     //290pi/512
   m_sin[291]  =  16'b1100000010000001;     //291pi/512
   m_cos[291]  =  16'b1111011111111110;     //291pi/512
   m_sin[292]  =  16'b1100000010001101;     //292pi/512
   m_cos[292]  =  16'b1111011110011111;     //292pi/512
   m_sin[293]  =  16'b1100000010011010;     //293pi/512
   m_cos[293]  =  16'b1111011101000000;     //293pi/512
   m_sin[294]  =  16'b1100000010100111;     //294pi/512
   m_cos[294]  =  16'b1111011011100010;     //294pi/512
   m_sin[295]  =  16'b1100000010110101;     //295pi/512
   m_cos[295]  =  16'b1111011010000011;     //295pi/512
   m_sin[296]  =  16'b1100000011000011;     //296pi/512
   m_cos[296]  =  16'b1111011000100101;     //296pi/512
   m_sin[297]  =  16'b1100000011010010;     //297pi/512
   m_cos[297]  =  16'b1111010111000110;     //297pi/512
   m_sin[298]  =  16'b1100000011100010;     //298pi/512
   m_cos[298]  =  16'b1111010101101000;     //298pi/512
   m_sin[299]  =  16'b1100000011110010;     //299pi/512
   m_cos[299]  =  16'b1111010100001010;     //299pi/512
   m_sin[300]  =  16'b1100000100000011;     //300pi/512
   m_cos[300]  =  16'b1111010010101100;     //300pi/512
   m_sin[301]  =  16'b1100000100010100;     //301pi/512
   m_cos[301]  =  16'b1111010001001110;     //301pi/512
   m_sin[302]  =  16'b1100000100100110;     //302pi/512
   m_cos[302]  =  16'b1111001111110000;     //302pi/512
   m_sin[303]  =  16'b1100000100111000;     //303pi/512
   m_cos[303]  =  16'b1111001110010010;     //303pi/512
   m_sin[304]  =  16'b1100000101001011;     //304pi/512
   m_cos[304]  =  16'b1111001100110101;     //304pi/512
   m_sin[305]  =  16'b1100000101011110;     //305pi/512
   m_cos[305]  =  16'b1111001011010111;     //305pi/512
   m_sin[306]  =  16'b1100000101110010;     //306pi/512
   m_cos[306]  =  16'b1111001001111010;     //306pi/512
   m_sin[307]  =  16'b1100000110000110;     //307pi/512
   m_cos[307]  =  16'b1111001000011101;     //307pi/512
   m_sin[308]  =  16'b1100000110011011;     //308pi/512
   m_cos[308]  =  16'b1111000110111111;     //308pi/512
   m_sin[309]  =  16'b1100000110110001;     //309pi/512
   m_cos[309]  =  16'b1111000101100010;     //309pi/512
   m_sin[310]  =  16'b1100000111000111;     //310pi/512
   m_cos[310]  =  16'b1111000100000101;     //310pi/512
   m_sin[311]  =  16'b1100000111011110;     //311pi/512
   m_cos[311]  =  16'b1111000010101001;     //311pi/512
   m_sin[312]  =  16'b1100000111110101;     //312pi/512
   m_cos[312]  =  16'b1111000001001100;     //312pi/512
   m_sin[313]  =  16'b1100001000001101;     //313pi/512
   m_cos[313]  =  16'b1110111111110000;     //313pi/512
   m_sin[314]  =  16'b1100001000100101;     //314pi/512
   m_cos[314]  =  16'b1110111110010011;     //314pi/512
   m_sin[315]  =  16'b1100001000111110;     //315pi/512
   m_cos[315]  =  16'b1110111100110111;     //315pi/512
   m_sin[316]  =  16'b1100001001010111;     //316pi/512
   m_cos[316]  =  16'b1110111011011011;     //316pi/512
   m_sin[317]  =  16'b1100001001110001;     //317pi/512
   m_cos[317]  =  16'b1110111001111111;     //317pi/512
   m_sin[318]  =  16'b1100001010001011;     //318pi/512
   m_cos[318]  =  16'b1110111000100011;     //318pi/512
   m_sin[319]  =  16'b1100001010100110;     //319pi/512
   m_cos[319]  =  16'b1110110111000111;     //319pi/512
   m_sin[320]  =  16'b1100001011000001;     //320pi/512
   m_cos[320]  =  16'b1110110101101100;     //320pi/512
   m_sin[321]  =  16'b1100001011011101;     //321pi/512
   m_cos[321]  =  16'b1110110100010001;     //321pi/512
   m_sin[322]  =  16'b1100001011111010;     //322pi/512
   m_cos[322]  =  16'b1110110010110110;     //322pi/512
   m_sin[323]  =  16'b1100001100010111;     //323pi/512
   m_cos[323]  =  16'b1110110001011011;     //323pi/512
   m_sin[324]  =  16'b1100001100110101;     //324pi/512
   m_cos[324]  =  16'b1110110000000000;     //324pi/512
   m_sin[325]  =  16'b1100001101010011;     //325pi/512
   m_cos[325]  =  16'b1110101110100101;     //325pi/512
   m_sin[326]  =  16'b1100001101110001;     //326pi/512
   m_cos[326]  =  16'b1110101101001011;     //326pi/512
   m_sin[327]  =  16'b1100001110010001;     //327pi/512
   m_cos[327]  =  16'b1110101011110000;     //327pi/512
   m_sin[328]  =  16'b1100001110110000;     //328pi/512
   m_cos[328]  =  16'b1110101010010110;     //328pi/512
   m_sin[329]  =  16'b1100001111010000;     //329pi/512
   m_cos[329]  =  16'b1110101000111100;     //329pi/512
   m_sin[330]  =  16'b1100001111110001;     //330pi/512
   m_cos[330]  =  16'b1110100111100011;     //330pi/512
   m_sin[331]  =  16'b1100010000010010;     //331pi/512
   m_cos[331]  =  16'b1110100110001001;     //331pi/512
   m_sin[332]  =  16'b1100010000110100;     //332pi/512
   m_cos[332]  =  16'b1110100100110000;     //332pi/512
   m_sin[333]  =  16'b1100010001010111;     //333pi/512
   m_cos[333]  =  16'b1110100011010111;     //333pi/512
   m_sin[334]  =  16'b1100010001111001;     //334pi/512
   m_cos[334]  =  16'b1110100001111110;     //334pi/512
   m_sin[335]  =  16'b1100010010011101;     //335pi/512
   m_cos[335]  =  16'b1110100000100101;     //335pi/512
   m_sin[336]  =  16'b1100010011000001;     //336pi/512
   m_cos[336]  =  16'b1110011111001100;     //336pi/512
   m_sin[337]  =  16'b1100010011100101;     //337pi/512
   m_cos[337]  =  16'b1110011101110100;     //337pi/512
   m_sin[338]  =  16'b1100010100001010;     //338pi/512
   m_cos[338]  =  16'b1110011100011100;     //338pi/512
   m_sin[339]  =  16'b1100010100101111;     //339pi/512
   m_cos[339]  =  16'b1110011011000100;     //339pi/512
   m_sin[340]  =  16'b1100010101010101;     //340pi/512
   m_cos[340]  =  16'b1110011001101101;     //340pi/512
   m_sin[341]  =  16'b1100010101111100;     //341pi/512
   m_cos[341]  =  16'b1110011000010101;     //341pi/512
   m_sin[342]  =  16'b1100010110100010;     //342pi/512
   m_cos[342]  =  16'b1110010110111110;     //342pi/512
   m_sin[343]  =  16'b1100010111001010;     //343pi/512
   m_cos[343]  =  16'b1110010101100111;     //343pi/512
   m_sin[344]  =  16'b1100010111110010;     //344pi/512
   m_cos[344]  =  16'b1110010100010000;     //344pi/512
   m_sin[345]  =  16'b1100011000011010;     //345pi/512
   m_cos[345]  =  16'b1110010010111010;     //345pi/512
   m_sin[346]  =  16'b1100011001000011;     //346pi/512
   m_cos[346]  =  16'b1110010001100011;     //346pi/512
   m_sin[347]  =  16'b1100011001101101;     //347pi/512
   m_cos[347]  =  16'b1110010000001101;     //347pi/512
   m_sin[348]  =  16'b1100011010010111;     //348pi/512
   m_cos[348]  =  16'b1110001110111000;     //348pi/512
   m_sin[349]  =  16'b1100011011000001;     //349pi/512
   m_cos[349]  =  16'b1110001101100010;     //349pi/512
   m_sin[350]  =  16'b1100011011101100;     //350pi/512
   m_cos[350]  =  16'b1110001100001101;     //350pi/512
   m_sin[351]  =  16'b1100011100011000;     //351pi/512
   m_cos[351]  =  16'b1110001010111000;     //351pi/512
   m_sin[352]  =  16'b1100011101000011;     //352pi/512
   m_cos[352]  =  16'b1110001001100011;     //352pi/512
   m_sin[353]  =  16'b1100011101110000;     //353pi/512
   m_cos[353]  =  16'b1110001000001110;     //353pi/512
   m_sin[354]  =  16'b1100011110011101;     //354pi/512
   m_cos[354]  =  16'b1110000110111010;     //354pi/512
   m_sin[355]  =  16'b1100011111001010;     //355pi/512
   m_cos[355]  =  16'b1110000101100110;     //355pi/512
   m_sin[356]  =  16'b1100011111111000;     //356pi/512
   m_cos[356]  =  16'b1110000100010010;     //356pi/512
   m_sin[357]  =  16'b1100100000100111;     //357pi/512
   m_cos[357]  =  16'b1110000010111111;     //357pi/512
   m_sin[358]  =  16'b1100100001010101;     //358pi/512
   m_cos[358]  =  16'b1110000001101100;     //358pi/512
   m_sin[359]  =  16'b1100100010000101;     //359pi/512
   m_cos[359]  =  16'b1110000000011001;     //359pi/512
   m_sin[360]  =  16'b1100100010110101;     //360pi/512
   m_cos[360]  =  16'b1101111111000110;     //360pi/512
   m_sin[361]  =  16'b1100100011100101;     //361pi/512
   m_cos[361]  =  16'b1101111101110100;     //361pi/512
   m_sin[362]  =  16'b1100100100010110;     //362pi/512
   m_cos[362]  =  16'b1101111100100010;     //362pi/512
   m_sin[363]  =  16'b1100100101000111;     //363pi/512
   m_cos[363]  =  16'b1101111011010000;     //363pi/512
   m_sin[364]  =  16'b1100100101111001;     //364pi/512
   m_cos[364]  =  16'b1101111001111110;     //364pi/512
   m_sin[365]  =  16'b1100100110101011;     //365pi/512
   m_cos[365]  =  16'b1101111000101101;     //365pi/512
   m_sin[366]  =  16'b1100100111011110;     //366pi/512
   m_cos[366]  =  16'b1101110111011100;     //366pi/512
   m_sin[367]  =  16'b1100101000010001;     //367pi/512
   m_cos[367]  =  16'b1101110110001011;     //367pi/512
   m_sin[368]  =  16'b1100101001000101;     //368pi/512
   m_cos[368]  =  16'b1101110100111011;     //368pi/512
   m_sin[369]  =  16'b1100101001111001;     //369pi/512
   m_cos[369]  =  16'b1101110011101011;     //369pi/512
   m_sin[370]  =  16'b1100101010101101;     //370pi/512
   m_cos[370]  =  16'b1101110010011011;     //370pi/512
   m_sin[371]  =  16'b1100101011100010;     //371pi/512
   m_cos[371]  =  16'b1101110001001100;     //371pi/512
   m_sin[372]  =  16'b1100101100011000;     //372pi/512
   m_cos[372]  =  16'b1101101111111101;     //372pi/512
   m_sin[373]  =  16'b1100101101001110;     //373pi/512
   m_cos[373]  =  16'b1101101110101110;     //373pi/512
   m_sin[374]  =  16'b1100101110000100;     //374pi/512
   m_cos[374]  =  16'b1101101101100000;     //374pi/512
   m_sin[375]  =  16'b1100101110111011;     //375pi/512
   m_cos[375]  =  16'b1101101100010001;     //375pi/512
   m_sin[376]  =  16'b1100101111110011;     //376pi/512
   m_cos[376]  =  16'b1101101011000100;     //376pi/512
   m_sin[377]  =  16'b1100110000101010;     //377pi/512
   m_cos[377]  =  16'b1101101001110110;     //377pi/512
   m_sin[378]  =  16'b1100110001100011;     //378pi/512
   m_cos[378]  =  16'b1101101000101001;     //378pi/512
   m_sin[379]  =  16'b1100110010011011;     //379pi/512
   m_cos[379]  =  16'b1101100111011100;     //379pi/512
   m_sin[380]  =  16'b1100110011010100;     //380pi/512
   m_cos[380]  =  16'b1101100110001111;     //380pi/512
   m_sin[381]  =  16'b1100110100001110;     //381pi/512
   m_cos[381]  =  16'b1101100101000011;     //381pi/512
   m_sin[382]  =  16'b1100110101001000;     //382pi/512
   m_cos[382]  =  16'b1101100011110111;     //382pi/512
   m_sin[383]  =  16'b1100110110000010;     //383pi/512
   m_cos[383]  =  16'b1101100010101100;     //383pi/512
   m_sin[384]  =  16'b1100110110111101;     //384pi/512
   m_cos[384]  =  16'b1101100001100001;     //384pi/512
   m_sin[385]  =  16'b1100110111111001;     //385pi/512
   m_cos[385]  =  16'b1101100000010110;     //385pi/512
   m_sin[386]  =  16'b1100111000110100;     //386pi/512
   m_cos[386]  =  16'b1101011111001011;     //386pi/512
   m_sin[387]  =  16'b1100111001110001;     //387pi/512
   m_cos[387]  =  16'b1101011110000001;     //387pi/512
   m_sin[388]  =  16'b1100111010101101;     //388pi/512
   m_cos[388]  =  16'b1101011100111000;     //388pi/512
   m_sin[389]  =  16'b1100111011101010;     //389pi/512
   m_cos[389]  =  16'b1101011011101110;     //389pi/512
   m_sin[390]  =  16'b1100111100101000;     //390pi/512
   m_cos[390]  =  16'b1101011010100101;     //390pi/512
   m_sin[391]  =  16'b1100111101100110;     //391pi/512
   m_cos[391]  =  16'b1101011001011100;     //391pi/512
   m_sin[392]  =  16'b1100111110100100;     //392pi/512
   m_cos[392]  =  16'b1101011000010100;     //392pi/512
   m_sin[393]  =  16'b1100111111100011;     //393pi/512
   m_cos[393]  =  16'b1101010111001100;     //393pi/512
   m_sin[394]  =  16'b1101000000100010;     //394pi/512
   m_cos[394]  =  16'b1101010110000100;     //394pi/512
   m_sin[395]  =  16'b1101000001100010;     //395pi/512
   m_cos[395]  =  16'b1101010100111101;     //395pi/512
   m_sin[396]  =  16'b1101000010100010;     //396pi/512
   m_cos[396]  =  16'b1101010011110110;     //396pi/512
   m_sin[397]  =  16'b1101000011100010;     //397pi/512
   m_cos[397]  =  16'b1101010010110000;     //397pi/512
   m_sin[398]  =  16'b1101000100100011;     //398pi/512
   m_cos[398]  =  16'b1101010001101010;     //398pi/512
   m_sin[399]  =  16'b1101000101100100;     //399pi/512
   m_cos[399]  =  16'b1101010000100100;     //399pi/512
   m_sin[400]  =  16'b1101000110100110;     //400pi/512
   m_cos[400]  =  16'b1101001111011111;     //400pi/512
   m_sin[401]  =  16'b1101000111101000;     //401pi/512
   m_cos[401]  =  16'b1101001110011010;     //401pi/512
   m_sin[402]  =  16'b1101001000101010;     //402pi/512
   m_cos[402]  =  16'b1101001101010101;     //402pi/512
   m_sin[403]  =  16'b1101001001101101;     //403pi/512
   m_cos[403]  =  16'b1101001100010001;     //403pi/512
   m_sin[404]  =  16'b1101001010110001;     //404pi/512
   m_cos[404]  =  16'b1101001011001101;     //404pi/512
   m_sin[405]  =  16'b1101001011110100;     //405pi/512
   m_cos[405]  =  16'b1101001010001010;     //405pi/512
   m_sin[406]  =  16'b1101001100111000;     //406pi/512
   m_cos[406]  =  16'b1101001001000111;     //406pi/512
   m_sin[407]  =  16'b1101001101111101;     //407pi/512
   m_cos[407]  =  16'b1101001000000100;     //407pi/512
   m_sin[408]  =  16'b1101001111000001;     //408pi/512
   m_cos[408]  =  16'b1101000111000010;     //408pi/512
   m_sin[409]  =  16'b1101010000000111;     //409pi/512
   m_cos[409]  =  16'b1101000110000000;     //409pi/512
   m_sin[410]  =  16'b1101010001001100;     //410pi/512
   m_cos[410]  =  16'b1101000100111110;     //410pi/512
   m_sin[411]  =  16'b1101010010010010;     //411pi/512
   m_cos[411]  =  16'b1101000011111101;     //411pi/512
   m_sin[412]  =  16'b1101010011011001;     //412pi/512
   m_cos[412]  =  16'b1101000010111101;     //412pi/512
   m_sin[413]  =  16'b1101010100011111;     //413pi/512
   m_cos[413]  =  16'b1101000001111101;     //413pi/512
   m_sin[414]  =  16'b1101010101100110;     //414pi/512
   m_cos[414]  =  16'b1101000000111101;     //414pi/512
   m_sin[415]  =  16'b1101010110101110;     //415pi/512
   m_cos[415]  =  16'b1100111111111110;     //415pi/512
   m_sin[416]  =  16'b1101010111110110;     //416pi/512
   m_cos[416]  =  16'b1100111110111111;     //416pi/512
   m_sin[417]  =  16'b1101011000111110;     //417pi/512
   m_cos[417]  =  16'b1100111110000000;     //417pi/512
   m_sin[418]  =  16'b1101011010000110;     //418pi/512
   m_cos[418]  =  16'b1100111101000010;     //418pi/512
   m_sin[419]  =  16'b1101011011001111;     //419pi/512
   m_cos[419]  =  16'b1100111100000100;     //419pi/512
   m_sin[420]  =  16'b1101011100011001;     //420pi/512
   m_cos[420]  =  16'b1100111011000111;     //420pi/512
   m_sin[421]  =  16'b1101011101100010;     //421pi/512
   m_cos[421]  =  16'b1100111010001010;     //421pi/512
   m_sin[422]  =  16'b1101011110101100;     //422pi/512
   m_cos[422]  =  16'b1100111001001110;     //422pi/512
   m_sin[423]  =  16'b1101011111110111;     //423pi/512
   m_cos[423]  =  16'b1100111000010010;     //423pi/512
   m_sin[424]  =  16'b1101100001000001;     //424pi/512
   m_cos[424]  =  16'b1100110111010110;     //424pi/512
   m_sin[425]  =  16'b1101100010001100;     //425pi/512
   m_cos[425]  =  16'b1100110110011011;     //425pi/512
   m_sin[426]  =  16'b1101100011011000;     //426pi/512
   m_cos[426]  =  16'b1100110101100001;     //426pi/512
   m_sin[427]  =  16'b1101100100100011;     //427pi/512
   m_cos[427]  =  16'b1100110100100110;     //427pi/512
   m_sin[428]  =  16'b1101100101101111;     //428pi/512
   m_cos[428]  =  16'b1100110011101101;     //428pi/512
   m_sin[429]  =  16'b1101100110111100;     //429pi/512
   m_cos[429]  =  16'b1100110010110011;     //429pi/512
   m_sin[430]  =  16'b1101101000001000;     //430pi/512
   m_cos[430]  =  16'b1100110001111010;     //430pi/512
   m_sin[431]  =  16'b1101101001010110;     //431pi/512
   m_cos[431]  =  16'b1100110001000010;     //431pi/512
   m_sin[432]  =  16'b1101101010100011;     //432pi/512
   m_cos[432]  =  16'b1100110000001010;     //432pi/512
   m_sin[433]  =  16'b1101101011110001;     //433pi/512
   m_cos[433]  =  16'b1100101111010010;     //433pi/512
   m_sin[434]  =  16'b1101101100111111;     //434pi/512
   m_cos[434]  =  16'b1100101110011011;     //434pi/512
   m_sin[435]  =  16'b1101101110001101;     //435pi/512
   m_cos[435]  =  16'b1100101101100101;     //435pi/512
   m_sin[436]  =  16'b1101101111011100;     //436pi/512
   m_cos[436]  =  16'b1100101100101111;     //436pi/512
   m_sin[437]  =  16'b1101110000101011;     //437pi/512
   m_cos[437]  =  16'b1100101011111001;     //437pi/512
   m_sin[438]  =  16'b1101110001111010;     //438pi/512
   m_cos[438]  =  16'b1100101011000100;     //438pi/512
   m_sin[439]  =  16'b1101110011001001;     //439pi/512
   m_cos[439]  =  16'b1100101010001111;     //439pi/512
   m_sin[440]  =  16'b1101110100011001;     //440pi/512
   m_cos[440]  =  16'b1100101001011011;     //440pi/512
   m_sin[441]  =  16'b1101110101101010;     //441pi/512
   m_cos[441]  =  16'b1100101000100111;     //441pi/512
   m_sin[442]  =  16'b1101110110111010;     //442pi/512
   m_cos[442]  =  16'b1100100111110011;     //442pi/512
   m_sin[443]  =  16'b1101111000001011;     //443pi/512
   m_cos[443]  =  16'b1100100111000000;     //443pi/512
   m_sin[444]  =  16'b1101111001011100;     //444pi/512
   m_cos[444]  =  16'b1100100110001110;     //444pi/512
   m_sin[445]  =  16'b1101111010101101;     //445pi/512
   m_cos[445]  =  16'b1100100101011100;     //445pi/512
   m_sin[446]  =  16'b1101111011111111;     //446pi/512
   m_cos[446]  =  16'b1100100100101011;     //446pi/512
   m_sin[447]  =  16'b1101111101010001;     //447pi/512
   m_cos[447]  =  16'b1100100011111001;     //447pi/512
   m_sin[448]  =  16'b1101111110100011;     //448pi/512
   m_cos[448]  =  16'b1100100011001001;     //448pi/512
   m_sin[449]  =  16'b1101111111110110;     //449pi/512
   m_cos[449]  =  16'b1100100010011001;     //449pi/512
   m_sin[450]  =  16'b1110000001001001;     //450pi/512
   m_cos[450]  =  16'b1100100001101001;     //450pi/512
   m_sin[451]  =  16'b1110000010011100;     //451pi/512
   m_cos[451]  =  16'b1100100000111010;     //451pi/512
   m_sin[452]  =  16'b1110000011101111;     //452pi/512
   m_cos[452]  =  16'b1100100000001100;     //452pi/512
   m_sin[453]  =  16'b1110000101000011;     //453pi/512
   m_cos[453]  =  16'b1100011111011110;     //453pi/512
   m_sin[454]  =  16'b1110000110010111;     //454pi/512
   m_cos[454]  =  16'b1100011110110000;     //454pi/512
   m_sin[455]  =  16'b1110000111101011;     //455pi/512
   m_cos[455]  =  16'b1100011110000011;     //455pi/512
   m_sin[456]  =  16'b1110001000111111;     //456pi/512
   m_cos[456]  =  16'b1100011101010110;     //456pi/512
   m_sin[457]  =  16'b1110001010010100;     //457pi/512
   m_cos[457]  =  16'b1100011100101010;     //457pi/512
   m_sin[458]  =  16'b1110001011101001;     //458pi/512
   m_cos[458]  =  16'b1100011011111110;     //458pi/512
   m_sin[459]  =  16'b1110001100111110;     //459pi/512
   m_cos[459]  =  16'b1100011011010011;     //459pi/512
   m_sin[460]  =  16'b1110001110010100;     //460pi/512
   m_cos[460]  =  16'b1100011010101000;     //460pi/512
   m_sin[461]  =  16'b1110001111101001;     //461pi/512
   m_cos[461]  =  16'b1100011001111110;     //461pi/512
   m_sin[462]  =  16'b1110010000111111;     //462pi/512
   m_cos[462]  =  16'b1100011001010101;     //462pi/512
   m_sin[463]  =  16'b1110010010010101;     //463pi/512
   m_cos[463]  =  16'b1100011000101011;     //463pi/512
   m_sin[464]  =  16'b1110010011101100;     //464pi/512
   m_cos[464]  =  16'b1100011000000011;     //464pi/512
   m_sin[465]  =  16'b1110010101000010;     //465pi/512
   m_cos[465]  =  16'b1100010111011011;     //465pi/512
   m_sin[466]  =  16'b1110010110011001;     //466pi/512
   m_cos[466]  =  16'b1100010110110011;     //466pi/512
   m_sin[467]  =  16'b1110010111110000;     //467pi/512
   m_cos[467]  =  16'b1100010110001100;     //467pi/512
   m_sin[468]  =  16'b1110011001001000;     //468pi/512
   m_cos[468]  =  16'b1100010101100101;     //468pi/512
   m_sin[469]  =  16'b1110011010011111;     //469pi/512
   m_cos[469]  =  16'b1100010100111111;     //469pi/512
   m_sin[470]  =  16'b1110011011110111;     //470pi/512
   m_cos[470]  =  16'b1100010100011010;     //470pi/512
   m_sin[471]  =  16'b1110011101001111;     //471pi/512
   m_cos[471]  =  16'b1100010011110100;     //471pi/512
   m_sin[472]  =  16'b1110011110100111;     //472pi/512
   m_cos[472]  =  16'b1100010011010000;     //472pi/512
   m_sin[473]  =  16'b1110100000000000;     //473pi/512
   m_cos[473]  =  16'b1100010010101100;     //473pi/512
   m_sin[474]  =  16'b1110100001011000;     //474pi/512
   m_cos[474]  =  16'b1100010010001000;     //474pi/512
   m_sin[475]  =  16'b1110100010110001;     //475pi/512
   m_cos[475]  =  16'b1100010001100101;     //475pi/512
   m_sin[476]  =  16'b1110100100001010;     //476pi/512
   m_cos[476]  =  16'b1100010001000011;     //476pi/512
   m_sin[477]  =  16'b1110100101100011;     //477pi/512
   m_cos[477]  =  16'b1100010000100001;     //477pi/512
   m_sin[478]  =  16'b1110100110111101;     //478pi/512
   m_cos[478]  =  16'b1100001111111111;     //478pi/512
   m_sin[479]  =  16'b1110101000010111;     //479pi/512
   m_cos[479]  =  16'b1100001111011110;     //479pi/512
   m_sin[480]  =  16'b1110101001110000;     //480pi/512
   m_cos[480]  =  16'b1100001110111110;     //480pi/512
   m_sin[481]  =  16'b1110101011001010;     //481pi/512
   m_cos[481]  =  16'b1100001110011110;     //481pi/512
   m_sin[482]  =  16'b1110101100100101;     //482pi/512
   m_cos[482]  =  16'b1100001101111110;     //482pi/512
   m_sin[483]  =  16'b1110101101111111;     //483pi/512
   m_cos[483]  =  16'b1100001101100000;     //483pi/512
   m_sin[484]  =  16'b1110101111011010;     //484pi/512
   m_cos[484]  =  16'b1100001101000001;     //484pi/512
   m_sin[485]  =  16'b1110110000110100;     //485pi/512
   m_cos[485]  =  16'b1100001100100011;     //485pi/512
   m_sin[486]  =  16'b1110110010001111;     //486pi/512
   m_cos[486]  =  16'b1100001100000110;     //486pi/512
   m_sin[487]  =  16'b1110110011101010;     //487pi/512
   m_cos[487]  =  16'b1100001011101001;     //487pi/512
   m_sin[488]  =  16'b1110110101000110;     //488pi/512
   m_cos[488]  =  16'b1100001011001101;     //488pi/512
   m_sin[489]  =  16'b1110110110100001;     //489pi/512
   m_cos[489]  =  16'b1100001010110010;     //489pi/512
   m_sin[490]  =  16'b1110110111111100;     //490pi/512
   m_cos[490]  =  16'b1100001010010110;     //490pi/512
   m_sin[491]  =  16'b1110111001011000;     //491pi/512
   m_cos[491]  =  16'b1100001001111100;     //491pi/512
   m_sin[492]  =  16'b1110111010110100;     //492pi/512
   m_cos[492]  =  16'b1100001001100010;     //492pi/512
   m_sin[493]  =  16'b1110111100010000;     //493pi/512
   m_cos[493]  =  16'b1100001001001000;     //493pi/512
   m_sin[494]  =  16'b1110111101101100;     //494pi/512
   m_cos[494]  =  16'b1100001000101111;     //494pi/512
   m_sin[495]  =  16'b1110111111001001;     //495pi/512
   m_cos[495]  =  16'b1100001000010111;     //495pi/512
   m_sin[496]  =  16'b1111000000100101;     //496pi/512
   m_cos[496]  =  16'b1100000111111111;     //496pi/512
   m_sin[497]  =  16'b1111000010000010;     //497pi/512
   m_cos[497]  =  16'b1100000111100111;     //497pi/512
   m_sin[498]  =  16'b1111000011011110;     //498pi/512
   m_cos[498]  =  16'b1100000111010001;     //498pi/512
   m_sin[499]  =  16'b1111000100111011;     //499pi/512
   m_cos[499]  =  16'b1100000110111010;     //499pi/512
   m_sin[500]  =  16'b1111000110011000;     //500pi/512
   m_cos[500]  =  16'b1100000110100100;     //500pi/512
   m_sin[501]  =  16'b1111000111110101;     //501pi/512
   m_cos[501]  =  16'b1100000110001111;     //501pi/512
   m_sin[502]  =  16'b1111001001010011;     //502pi/512
   m_cos[502]  =  16'b1100000101111011;     //502pi/512
   m_sin[503]  =  16'b1111001010110000;     //503pi/512
   m_cos[503]  =  16'b1100000101100110;     //503pi/512
   m_sin[504]  =  16'b1111001100001101;     //504pi/512
   m_cos[504]  =  16'b1100000101010011;     //504pi/512
   m_sin[505]  =  16'b1111001101101011;     //505pi/512
   m_cos[505]  =  16'b1100000101000000;     //505pi/512
   m_sin[506]  =  16'b1111001111001001;     //506pi/512
   m_cos[506]  =  16'b1100000100101101;     //506pi/512
   m_sin[507]  =  16'b1111010000100110;     //507pi/512
   m_cos[507]  =  16'b1100000100011011;     //507pi/512
   m_sin[508]  =  16'b1111010010000100;     //508pi/512
   m_cos[508]  =  16'b1100000100001010;     //508pi/512
   m_sin[509]  =  16'b1111010011100010;     //509pi/512
   m_cos[509]  =  16'b1100000011111001;     //509pi/512
   m_sin[510]  =  16'b1111010101000000;     //510pi/512
   m_cos[510]  =  16'b1100000011101001;     //510pi/512
   m_sin[511]  =  16'b1111010110011111;     //511pi/512
   m_cos[511]  =  16'b1100000011011001;     //511pi/512
end
endmodule
