module  M_TWIDLE_14_B_0_15_v #(parameter SIZE =10, word_length_tw = 14) (
    input            clk,
    input            en_rd, 
    input   [10:0]   rd_ptr_angle,
    input            en_modf, 

    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );


reg signed [word_length_tw-1:0]  cos  [511:0];
reg signed [word_length_tw-1:0]  sin  [511:0];

reg signed [word_length_tw-1:0]  m_cos  [511:0];
reg signed [word_length_tw-1:0]  m_sin  [511:0];

reg signed [word_length_tw-1:0]  cos_temp;
reg signed [word_length_tw-1:0]  sin_temp;

reg signed [word_length_tw-1:0]  m_cos_temp;
reg signed [word_length_tw-1:0]  m_sin_temp;


//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & ~ en_modf ) begin
                  cos_temp           <= cos   [rd_ptr_angle];
                  sin_temp           <= sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & en_modf ) begin
                  m_cos_temp           <= m_cos   [rd_ptr_angle];
                  m_sin_temp           <= m_sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(*) begin 
             if (en_modf ) begin
                  cos_data           <= m_cos_temp;
                  sin_data           <= m_sin_temp;
             end else begin
                  cos_data           <= cos_temp;
                  sin_data           <= sin_temp;
             end
        end
//----------------------------------------------------------------------------------------
initial begin
   sin[0]  =  14'b00000000000000;     //0pi/512
   cos[0]  =  14'b01000000000000;     //0pi/512
   sin[1]  =  14'b11111111100111;     //1pi/512
   cos[1]  =  14'b00111111111111;     //1pi/512
   sin[2]  =  14'b11111111001110;     //2pi/512
   cos[2]  =  14'b00111111111111;     //2pi/512
   sin[3]  =  14'b11111110110101;     //3pi/512
   cos[3]  =  14'b00111111111111;     //3pi/512
   sin[4]  =  14'b11111110011011;     //4pi/512
   cos[4]  =  14'b00111111111110;     //4pi/512
   sin[5]  =  14'b11111110000010;     //5pi/512
   cos[5]  =  14'b00111111111110;     //5pi/512
   sin[6]  =  14'b11111101101001;     //6pi/512
   cos[6]  =  14'b00111111111101;     //6pi/512
   sin[7]  =  14'b11111101010000;     //7pi/512
   cos[7]  =  14'b00111111111100;     //7pi/512
   sin[8]  =  14'b11111100110111;     //8pi/512
   cos[8]  =  14'b00111111111011;     //8pi/512
   sin[9]  =  14'b11111100011110;     //9pi/512
   cos[9]  =  14'b00111111111001;     //9pi/512
   sin[10]  =  14'b11111100000101;     //10pi/512
   cos[10]  =  14'b00111111111000;     //10pi/512
   sin[11]  =  14'b11111011101100;     //11pi/512
   cos[11]  =  14'b00111111110110;     //11pi/512
   sin[12]  =  14'b11111011010011;     //12pi/512
   cos[12]  =  14'b00111111110100;     //12pi/512
   sin[13]  =  14'b11111010111010;     //13pi/512
   cos[13]  =  14'b00111111110010;     //13pi/512
   sin[14]  =  14'b11111010100001;     //14pi/512
   cos[14]  =  14'b00111111110000;     //14pi/512
   sin[15]  =  14'b11111010001000;     //15pi/512
   cos[15]  =  14'b00111111101110;     //15pi/512
   sin[16]  =  14'b11111001101111;     //16pi/512
   cos[16]  =  14'b00111111101100;     //16pi/512
   sin[17]  =  14'b11111001010110;     //17pi/512
   cos[17]  =  14'b00111111101001;     //17pi/512
   sin[18]  =  14'b11111000111101;     //18pi/512
   cos[18]  =  14'b00111111100111;     //18pi/512
   sin[19]  =  14'b11111000100100;     //19pi/512
   cos[19]  =  14'b00111111100100;     //19pi/512
   sin[20]  =  14'b11111000001011;     //20pi/512
   cos[20]  =  14'b00111111100001;     //20pi/512
   sin[21]  =  14'b11110111110010;     //21pi/512
   cos[21]  =  14'b00111111011110;     //21pi/512
   sin[22]  =  14'b11110111011001;     //22pi/512
   cos[22]  =  14'b00111111011010;     //22pi/512
   sin[23]  =  14'b11110111000000;     //23pi/512
   cos[23]  =  14'b00111111010111;     //23pi/512
   sin[24]  =  14'b11110110100111;     //24pi/512
   cos[24]  =  14'b00111111010011;     //24pi/512
   sin[25]  =  14'b11110110001110;     //25pi/512
   cos[25]  =  14'b00111111001111;     //25pi/512
   sin[26]  =  14'b11110101110101;     //26pi/512
   cos[26]  =  14'b00111111001011;     //26pi/512
   sin[27]  =  14'b11110101011101;     //27pi/512
   cos[27]  =  14'b00111111000111;     //27pi/512
   sin[28]  =  14'b11110101000100;     //28pi/512
   cos[28]  =  14'b00111111000011;     //28pi/512
   sin[29]  =  14'b11110100101011;     //29pi/512
   cos[29]  =  14'b00111110111111;     //29pi/512
   sin[30]  =  14'b11110100010010;     //30pi/512
   cos[30]  =  14'b00111110111010;     //30pi/512
   sin[31]  =  14'b11110011111010;     //31pi/512
   cos[31]  =  14'b00111110110110;     //31pi/512
   sin[32]  =  14'b11110011100001;     //32pi/512
   cos[32]  =  14'b00111110110001;     //32pi/512
   sin[33]  =  14'b11110011001000;     //33pi/512
   cos[33]  =  14'b00111110101100;     //33pi/512
   sin[34]  =  14'b11110010110000;     //34pi/512
   cos[34]  =  14'b00111110100111;     //34pi/512
   sin[35]  =  14'b11110010010111;     //35pi/512
   cos[35]  =  14'b00111110100001;     //35pi/512
   sin[36]  =  14'b11110001111111;     //36pi/512
   cos[36]  =  14'b00111110011100;     //36pi/512
   sin[37]  =  14'b11110001100110;     //37pi/512
   cos[37]  =  14'b00111110010110;     //37pi/512
   sin[38]  =  14'b11110001001110;     //38pi/512
   cos[38]  =  14'b00111110010001;     //38pi/512
   sin[39]  =  14'b11110000110101;     //39pi/512
   cos[39]  =  14'b00111110001011;     //39pi/512
   sin[40]  =  14'b11110000011101;     //40pi/512
   cos[40]  =  14'b00111110000101;     //40pi/512
   sin[41]  =  14'b11110000000100;     //41pi/512
   cos[41]  =  14'b00111101111111;     //41pi/512
   sin[42]  =  14'b11101111101100;     //42pi/512
   cos[42]  =  14'b00111101111000;     //42pi/512
   sin[43]  =  14'b11101111010100;     //43pi/512
   cos[43]  =  14'b00111101110010;     //43pi/512
   sin[44]  =  14'b11101110111100;     //44pi/512
   cos[44]  =  14'b00111101101011;     //44pi/512
   sin[45]  =  14'b11101110100011;     //45pi/512
   cos[45]  =  14'b00111101100100;     //45pi/512
   sin[46]  =  14'b11101110001011;     //46pi/512
   cos[46]  =  14'b00111101011101;     //46pi/512
   sin[47]  =  14'b11101101110011;     //47pi/512
   cos[47]  =  14'b00111101010110;     //47pi/512
   sin[48]  =  14'b11101101011011;     //48pi/512
   cos[48]  =  14'b00111101001111;     //48pi/512
   sin[49]  =  14'b11101101000011;     //49pi/512
   cos[49]  =  14'b00111101001000;     //49pi/512
   sin[50]  =  14'b11101100101011;     //50pi/512
   cos[50]  =  14'b00111101000000;     //50pi/512
   sin[51]  =  14'b11101100010011;     //51pi/512
   cos[51]  =  14'b00111100111001;     //51pi/512
   sin[52]  =  14'b11101011111011;     //52pi/512
   cos[52]  =  14'b00111100110001;     //52pi/512
   sin[53]  =  14'b11101011100011;     //53pi/512
   cos[53]  =  14'b00111100101001;     //53pi/512
   sin[54]  =  14'b11101011001100;     //54pi/512
   cos[54]  =  14'b00111100100001;     //54pi/512
   sin[55]  =  14'b11101010110100;     //55pi/512
   cos[55]  =  14'b00111100011000;     //55pi/512
   sin[56]  =  14'b11101010011100;     //56pi/512
   cos[56]  =  14'b00111100010000;     //56pi/512
   sin[57]  =  14'b11101010000100;     //57pi/512
   cos[57]  =  14'b00111100001000;     //57pi/512
   sin[58]  =  14'b11101001101101;     //58pi/512
   cos[58]  =  14'b00111011111111;     //58pi/512
   sin[59]  =  14'b11101001010101;     //59pi/512
   cos[59]  =  14'b00111011110110;     //59pi/512
   sin[60]  =  14'b11101000111110;     //60pi/512
   cos[60]  =  14'b00111011101101;     //60pi/512
   sin[61]  =  14'b11101000100110;     //61pi/512
   cos[61]  =  14'b00111011100100;     //61pi/512
   sin[62]  =  14'b11101000001111;     //62pi/512
   cos[62]  =  14'b00111011011011;     //62pi/512
   sin[63]  =  14'b11100111111000;     //63pi/512
   cos[63]  =  14'b00111011010001;     //63pi/512
   sin[64]  =  14'b11100111100001;     //64pi/512
   cos[64]  =  14'b00111011001000;     //64pi/512
   sin[65]  =  14'b11100111001001;     //65pi/512
   cos[65]  =  14'b00111010111110;     //65pi/512
   sin[66]  =  14'b11100110110010;     //66pi/512
   cos[66]  =  14'b00111010110100;     //66pi/512
   sin[67]  =  14'b11100110011011;     //67pi/512
   cos[67]  =  14'b00111010101010;     //67pi/512
   sin[68]  =  14'b11100110000100;     //68pi/512
   cos[68]  =  14'b00111010100000;     //68pi/512
   sin[69]  =  14'b11100101101101;     //69pi/512
   cos[69]  =  14'b00111010010110;     //69pi/512
   sin[70]  =  14'b11100101010110;     //70pi/512
   cos[70]  =  14'b00111010001011;     //70pi/512
   sin[71]  =  14'b11100100111111;     //71pi/512
   cos[71]  =  14'b00111010000001;     //71pi/512
   sin[72]  =  14'b11100100101001;     //72pi/512
   cos[72]  =  14'b00111001110110;     //72pi/512
   sin[73]  =  14'b11100100010010;     //73pi/512
   cos[73]  =  14'b00111001101011;     //73pi/512
   sin[74]  =  14'b11100011111011;     //74pi/512
   cos[74]  =  14'b00111001100000;     //74pi/512
   sin[75]  =  14'b11100011100101;     //75pi/512
   cos[75]  =  14'b00111001010101;     //75pi/512
   sin[76]  =  14'b11100011001110;     //76pi/512
   cos[76]  =  14'b00111001001010;     //76pi/512
   sin[77]  =  14'b11100010111000;     //77pi/512
   cos[77]  =  14'b00111000111111;     //77pi/512
   sin[78]  =  14'b11100010100010;     //78pi/512
   cos[78]  =  14'b00111000110011;     //78pi/512
   sin[79]  =  14'b11100010001011;     //79pi/512
   cos[79]  =  14'b00111000101000;     //79pi/512
   sin[80]  =  14'b11100001110101;     //80pi/512
   cos[80]  =  14'b00111000011100;     //80pi/512
   sin[81]  =  14'b11100001011111;     //81pi/512
   cos[81]  =  14'b00111000010000;     //81pi/512
   sin[82]  =  14'b11100001001001;     //82pi/512
   cos[82]  =  14'b00111000000100;     //82pi/512
   sin[83]  =  14'b11100000110011;     //83pi/512
   cos[83]  =  14'b00110111111000;     //83pi/512
   sin[84]  =  14'b11100000011101;     //84pi/512
   cos[84]  =  14'b00110111101011;     //84pi/512
   sin[85]  =  14'b11100000000111;     //85pi/512
   cos[85]  =  14'b00110111011111;     //85pi/512
   sin[86]  =  14'b11011111110010;     //86pi/512
   cos[86]  =  14'b00110111010010;     //86pi/512
   sin[87]  =  14'b11011111011100;     //87pi/512
   cos[87]  =  14'b00110111000110;     //87pi/512
   sin[88]  =  14'b11011111000110;     //88pi/512
   cos[88]  =  14'b00110110111001;     //88pi/512
   sin[89]  =  14'b11011110110001;     //89pi/512
   cos[89]  =  14'b00110110101100;     //89pi/512
   sin[90]  =  14'b11011110011011;     //90pi/512
   cos[90]  =  14'b00110110011111;     //90pi/512
   sin[91]  =  14'b11011110000110;     //91pi/512
   cos[91]  =  14'b00110110010001;     //91pi/512
   sin[92]  =  14'b11011101110001;     //92pi/512
   cos[92]  =  14'b00110110000100;     //92pi/512
   sin[93]  =  14'b11011101011011;     //93pi/512
   cos[93]  =  14'b00110101110111;     //93pi/512
   sin[94]  =  14'b11011101000110;     //94pi/512
   cos[94]  =  14'b00110101101001;     //94pi/512
   sin[95]  =  14'b11011100110001;     //95pi/512
   cos[95]  =  14'b00110101011011;     //95pi/512
   sin[96]  =  14'b11011100011100;     //96pi/512
   cos[96]  =  14'b00110101001101;     //96pi/512
   sin[97]  =  14'b11011100001000;     //97pi/512
   cos[97]  =  14'b00110100111111;     //97pi/512
   sin[98]  =  14'b11011011110011;     //98pi/512
   cos[98]  =  14'b00110100110001;     //98pi/512
   sin[99]  =  14'b11011011011110;     //99pi/512
   cos[99]  =  14'b00110100100011;     //99pi/512
   sin[100]  =  14'b11011011001001;     //100pi/512
   cos[100]  =  14'b00110100010100;     //100pi/512
   sin[101]  =  14'b11011010110101;     //101pi/512
   cos[101]  =  14'b00110100000110;     //101pi/512
   sin[102]  =  14'b11011010100001;     //102pi/512
   cos[102]  =  14'b00110011110111;     //102pi/512
   sin[103]  =  14'b11011010001100;     //103pi/512
   cos[103]  =  14'b00110011101000;     //103pi/512
   sin[104]  =  14'b11011001111000;     //104pi/512
   cos[104]  =  14'b00110011011001;     //104pi/512
   sin[105]  =  14'b11011001100100;     //105pi/512
   cos[105]  =  14'b00110011001010;     //105pi/512
   sin[106]  =  14'b11011001010000;     //106pi/512
   cos[106]  =  14'b00110010111011;     //106pi/512
   sin[107]  =  14'b11011000111100;     //107pi/512
   cos[107]  =  14'b00110010101100;     //107pi/512
   sin[108]  =  14'b11011000101000;     //108pi/512
   cos[108]  =  14'b00110010011101;     //108pi/512
   sin[109]  =  14'b11011000010100;     //109pi/512
   cos[109]  =  14'b00110010001101;     //109pi/512
   sin[110]  =  14'b11011000000001;     //110pi/512
   cos[110]  =  14'b00110001111101;     //110pi/512
   sin[111]  =  14'b11010111101101;     //111pi/512
   cos[111]  =  14'b00110001101110;     //111pi/512
   sin[112]  =  14'b11010111011010;     //112pi/512
   cos[112]  =  14'b00110001011110;     //112pi/512
   sin[113]  =  14'b11010111000110;     //113pi/512
   cos[113]  =  14'b00110001001110;     //113pi/512
   sin[114]  =  14'b11010110110011;     //114pi/512
   cos[114]  =  14'b00110000111110;     //114pi/512
   sin[115]  =  14'b11010110100000;     //115pi/512
   cos[115]  =  14'b00110000101101;     //115pi/512
   sin[116]  =  14'b11010110001101;     //116pi/512
   cos[116]  =  14'b00110000011101;     //116pi/512
   sin[117]  =  14'b11010101111010;     //117pi/512
   cos[117]  =  14'b00110000001101;     //117pi/512
   sin[118]  =  14'b11010101100111;     //118pi/512
   cos[118]  =  14'b00101111111100;     //118pi/512
   sin[119]  =  14'b11010101010100;     //119pi/512
   cos[119]  =  14'b00101111101011;     //119pi/512
   sin[120]  =  14'b11010101000001;     //120pi/512
   cos[120]  =  14'b00101111011010;     //120pi/512
   sin[121]  =  14'b11010100101111;     //121pi/512
   cos[121]  =  14'b00101111001010;     //121pi/512
   sin[122]  =  14'b11010100011100;     //122pi/512
   cos[122]  =  14'b00101110111000;     //122pi/512
   sin[123]  =  14'b11010100001010;     //123pi/512
   cos[123]  =  14'b00101110100111;     //123pi/512
   sin[124]  =  14'b11010011111000;     //124pi/512
   cos[124]  =  14'b00101110010110;     //124pi/512
   sin[125]  =  14'b11010011100101;     //125pi/512
   cos[125]  =  14'b00101110000101;     //125pi/512
   sin[126]  =  14'b11010011010011;     //126pi/512
   cos[126]  =  14'b00101101110011;     //126pi/512
   sin[127]  =  14'b11010011000010;     //127pi/512
   cos[127]  =  14'b00101101100010;     //127pi/512
   sin[128]  =  14'b11010010110000;     //128pi/512
   cos[128]  =  14'b00101101010000;     //128pi/512
   sin[129]  =  14'b11010010011110;     //129pi/512
   cos[129]  =  14'b00101100111110;     //129pi/512
   sin[130]  =  14'b11010010001100;     //130pi/512
   cos[130]  =  14'b00101100101100;     //130pi/512
   sin[131]  =  14'b11010001111011;     //131pi/512
   cos[131]  =  14'b00101100011010;     //131pi/512
   sin[132]  =  14'b11010001101001;     //132pi/512
   cos[132]  =  14'b00101100001000;     //132pi/512
   sin[133]  =  14'b11010001011000;     //133pi/512
   cos[133]  =  14'b00101011110110;     //133pi/512
   sin[134]  =  14'b11010001000111;     //134pi/512
   cos[134]  =  14'b00101011100011;     //134pi/512
   sin[135]  =  14'b11010000110110;     //135pi/512
   cos[135]  =  14'b00101011010001;     //135pi/512
   sin[136]  =  14'b11010000100101;     //136pi/512
   cos[136]  =  14'b00101010111110;     //136pi/512
   sin[137]  =  14'b11010000010100;     //137pi/512
   cos[137]  =  14'b00101010101100;     //137pi/512
   sin[138]  =  14'b11010000000100;     //138pi/512
   cos[138]  =  14'b00101010011001;     //138pi/512
   sin[139]  =  14'b11001111110011;     //139pi/512
   cos[139]  =  14'b00101010000110;     //139pi/512
   sin[140]  =  14'b11001111100010;     //140pi/512
   cos[140]  =  14'b00101001110011;     //140pi/512
   sin[141]  =  14'b11001111010010;     //141pi/512
   cos[141]  =  14'b00101001100000;     //141pi/512
   sin[142]  =  14'b11001111000010;     //142pi/512
   cos[142]  =  14'b00101001001101;     //142pi/512
   sin[143]  =  14'b11001110110010;     //143pi/512
   cos[143]  =  14'b00101000111001;     //143pi/512
   sin[144]  =  14'b11001110100010;     //144pi/512
   cos[144]  =  14'b00101000100110;     //144pi/512
   sin[145]  =  14'b11001110010010;     //145pi/512
   cos[145]  =  14'b00101000010010;     //145pi/512
   sin[146]  =  14'b11001110000010;     //146pi/512
   cos[146]  =  14'b00100111111111;     //146pi/512
   sin[147]  =  14'b11001101110010;     //147pi/512
   cos[147]  =  14'b00100111101011;     //147pi/512
   sin[148]  =  14'b11001101100011;     //148pi/512
   cos[148]  =  14'b00100111010111;     //148pi/512
   sin[149]  =  14'b11001101010100;     //149pi/512
   cos[149]  =  14'b00100111000100;     //149pi/512
   sin[150]  =  14'b11001101000100;     //150pi/512
   cos[150]  =  14'b00100110110000;     //150pi/512
   sin[151]  =  14'b11001100110101;     //151pi/512
   cos[151]  =  14'b00100110011100;     //151pi/512
   sin[152]  =  14'b11001100100110;     //152pi/512
   cos[152]  =  14'b00100110000111;     //152pi/512
   sin[153]  =  14'b11001100010111;     //153pi/512
   cos[153]  =  14'b00100101110011;     //153pi/512
   sin[154]  =  14'b11001100001000;     //154pi/512
   cos[154]  =  14'b00100101011111;     //154pi/512
   sin[155]  =  14'b11001011111010;     //155pi/512
   cos[155]  =  14'b00100101001011;     //155pi/512
   sin[156]  =  14'b11001011101011;     //156pi/512
   cos[156]  =  14'b00100100110110;     //156pi/512
   sin[157]  =  14'b11001011011101;     //157pi/512
   cos[157]  =  14'b00100100100001;     //157pi/512
   sin[158]  =  14'b11001011001110;     //158pi/512
   cos[158]  =  14'b00100100001101;     //158pi/512
   sin[159]  =  14'b11001011000000;     //159pi/512
   cos[159]  =  14'b00100011111000;     //159pi/512
   sin[160]  =  14'b11001010110010;     //160pi/512
   cos[160]  =  14'b00100011100011;     //160pi/512
   sin[161]  =  14'b11001010100100;     //161pi/512
   cos[161]  =  14'b00100011001110;     //161pi/512
   sin[162]  =  14'b11001010010111;     //162pi/512
   cos[162]  =  14'b00100010111001;     //162pi/512
   sin[163]  =  14'b11001010001001;     //163pi/512
   cos[163]  =  14'b00100010100100;     //163pi/512
   sin[164]  =  14'b11001001111011;     //164pi/512
   cos[164]  =  14'b00100010001111;     //164pi/512
   sin[165]  =  14'b11001001101110;     //165pi/512
   cos[165]  =  14'b00100001111010;     //165pi/512
   sin[166]  =  14'b11001001100001;     //166pi/512
   cos[166]  =  14'b00100001100100;     //166pi/512
   sin[167]  =  14'b11001001010100;     //167pi/512
   cos[167]  =  14'b00100001001111;     //167pi/512
   sin[168]  =  14'b11001001000111;     //168pi/512
   cos[168]  =  14'b00100000111001;     //168pi/512
   sin[169]  =  14'b11001000111010;     //169pi/512
   cos[169]  =  14'b00100000100100;     //169pi/512
   sin[170]  =  14'b11001000101101;     //170pi/512
   cos[170]  =  14'b00100000001110;     //170pi/512
   sin[171]  =  14'b11001000100001;     //171pi/512
   cos[171]  =  14'b00011111111000;     //171pi/512
   sin[172]  =  14'b11001000010100;     //172pi/512
   cos[172]  =  14'b00011111100010;     //172pi/512
   sin[173]  =  14'b11001000001000;     //173pi/512
   cos[173]  =  14'b00011111001101;     //173pi/512
   sin[174]  =  14'b11000111111100;     //174pi/512
   cos[174]  =  14'b00011110110111;     //174pi/512
   sin[175]  =  14'b11000111110000;     //175pi/512
   cos[175]  =  14'b00011110100000;     //175pi/512
   sin[176]  =  14'b11000111100100;     //176pi/512
   cos[176]  =  14'b00011110001010;     //176pi/512
   sin[177]  =  14'b11000111011000;     //177pi/512
   cos[177]  =  14'b00011101110100;     //177pi/512
   sin[178]  =  14'b11000111001100;     //178pi/512
   cos[178]  =  14'b00011101011110;     //178pi/512
   sin[179]  =  14'b11000111000001;     //179pi/512
   cos[179]  =  14'b00011101001000;     //179pi/512
   sin[180]  =  14'b11000110110101;     //180pi/512
   cos[180]  =  14'b00011100110001;     //180pi/512
   sin[181]  =  14'b11000110101010;     //181pi/512
   cos[181]  =  14'b00011100011011;     //181pi/512
   sin[182]  =  14'b11000110011111;     //182pi/512
   cos[182]  =  14'b00011100000100;     //182pi/512
   sin[183]  =  14'b11000110010100;     //183pi/512
   cos[183]  =  14'b00011011101101;     //183pi/512
   sin[184]  =  14'b11000110001001;     //184pi/512
   cos[184]  =  14'b00011011010111;     //184pi/512
   sin[185]  =  14'b11000101111111;     //185pi/512
   cos[185]  =  14'b00011011000000;     //185pi/512
   sin[186]  =  14'b11000101110100;     //186pi/512
   cos[186]  =  14'b00011010101001;     //186pi/512
   sin[187]  =  14'b11000101101010;     //187pi/512
   cos[187]  =  14'b00011010010010;     //187pi/512
   sin[188]  =  14'b11000101011111;     //188pi/512
   cos[188]  =  14'b00011001111011;     //188pi/512
   sin[189]  =  14'b11000101010101;     //189pi/512
   cos[189]  =  14'b00011001100100;     //189pi/512
   sin[190]  =  14'b11000101001011;     //190pi/512
   cos[190]  =  14'b00011001001101;     //190pi/512
   sin[191]  =  14'b11000101000001;     //191pi/512
   cos[191]  =  14'b00011000110110;     //191pi/512
   sin[192]  =  14'b11000100111000;     //192pi/512
   cos[192]  =  14'b00011000011111;     //192pi/512
   sin[193]  =  14'b11000100101110;     //193pi/512
   cos[193]  =  14'b00011000001000;     //193pi/512
   sin[194]  =  14'b11000100100101;     //194pi/512
   cos[194]  =  14'b00010111110000;     //194pi/512
   sin[195]  =  14'b11000100011100;     //195pi/512
   cos[195]  =  14'b00010111011001;     //195pi/512
   sin[196]  =  14'b11000100010010;     //196pi/512
   cos[196]  =  14'b00010111000010;     //196pi/512
   sin[197]  =  14'b11000100001001;     //197pi/512
   cos[197]  =  14'b00010110101010;     //197pi/512
   sin[198]  =  14'b11000100000001;     //198pi/512
   cos[198]  =  14'b00010110010011;     //198pi/512
   sin[199]  =  14'b11000011111000;     //199pi/512
   cos[199]  =  14'b00010101111011;     //199pi/512
   sin[200]  =  14'b11000011101111;     //200pi/512
   cos[200]  =  14'b00010101100011;     //200pi/512
   sin[201]  =  14'b11000011100111;     //201pi/512
   cos[201]  =  14'b00010101001100;     //201pi/512
   sin[202]  =  14'b11000011011111;     //202pi/512
   cos[202]  =  14'b00010100110100;     //202pi/512
   sin[203]  =  14'b11000011010111;     //203pi/512
   cos[203]  =  14'b00010100011100;     //203pi/512
   sin[204]  =  14'b11000011001111;     //204pi/512
   cos[204]  =  14'b00010100000100;     //204pi/512
   sin[205]  =  14'b11000011000111;     //205pi/512
   cos[205]  =  14'b00010011101100;     //205pi/512
   sin[206]  =  14'b11000010111111;     //206pi/512
   cos[206]  =  14'b00010011010101;     //206pi/512
   sin[207]  =  14'b11000010111000;     //207pi/512
   cos[207]  =  14'b00010010111101;     //207pi/512
   sin[208]  =  14'b11000010110000;     //208pi/512
   cos[208]  =  14'b00010010100101;     //208pi/512
   sin[209]  =  14'b11000010101001;     //209pi/512
   cos[209]  =  14'b00010010001100;     //209pi/512
   sin[210]  =  14'b11000010100010;     //210pi/512
   cos[210]  =  14'b00010001110100;     //210pi/512
   sin[211]  =  14'b11000010011011;     //211pi/512
   cos[211]  =  14'b00010001011100;     //211pi/512
   sin[212]  =  14'b11000010010100;     //212pi/512
   cos[212]  =  14'b00010001000100;     //212pi/512
   sin[213]  =  14'b11000010001110;     //213pi/512
   cos[213]  =  14'b00010000101100;     //213pi/512
   sin[214]  =  14'b11000010000111;     //214pi/512
   cos[214]  =  14'b00010000010011;     //214pi/512
   sin[215]  =  14'b11000010000001;     //215pi/512
   cos[215]  =  14'b00001111111011;     //215pi/512
   sin[216]  =  14'b11000001111011;     //216pi/512
   cos[216]  =  14'b00001111100011;     //216pi/512
   sin[217]  =  14'b11000001110101;     //217pi/512
   cos[217]  =  14'b00001111001010;     //217pi/512
   sin[218]  =  14'b11000001101111;     //218pi/512
   cos[218]  =  14'b00001110110010;     //218pi/512
   sin[219]  =  14'b11000001101001;     //219pi/512
   cos[219]  =  14'b00001110011001;     //219pi/512
   sin[220]  =  14'b11000001100100;     //220pi/512
   cos[220]  =  14'b00001110000001;     //220pi/512
   sin[221]  =  14'b11000001011110;     //221pi/512
   cos[221]  =  14'b00001101101000;     //221pi/512
   sin[222]  =  14'b11000001011001;     //222pi/512
   cos[222]  =  14'b00001101010000;     //222pi/512
   sin[223]  =  14'b11000001010100;     //223pi/512
   cos[223]  =  14'b00001100110111;     //223pi/512
   sin[224]  =  14'b11000001001111;     //224pi/512
   cos[224]  =  14'b00001100011111;     //224pi/512
   sin[225]  =  14'b11000001001010;     //225pi/512
   cos[225]  =  14'b00001100000110;     //225pi/512
   sin[226]  =  14'b11000001000101;     //226pi/512
   cos[226]  =  14'b00001011101101;     //226pi/512
   sin[227]  =  14'b11000001000001;     //227pi/512
   cos[227]  =  14'b00001011010101;     //227pi/512
   sin[228]  =  14'b11000000111100;     //228pi/512
   cos[228]  =  14'b00001010111100;     //228pi/512
   sin[229]  =  14'b11000000111000;     //229pi/512
   cos[229]  =  14'b00001010100011;     //229pi/512
   sin[230]  =  14'b11000000110100;     //230pi/512
   cos[230]  =  14'b00001010001010;     //230pi/512
   sin[231]  =  14'b11000000110000;     //231pi/512
   cos[231]  =  14'b00001001110001;     //231pi/512
   sin[232]  =  14'b11000000101100;     //232pi/512
   cos[232]  =  14'b00001001011001;     //232pi/512
   sin[233]  =  14'b11000000101001;     //233pi/512
   cos[233]  =  14'b00001001000000;     //233pi/512
   sin[234]  =  14'b11000000100101;     //234pi/512
   cos[234]  =  14'b00001000100111;     //234pi/512
   sin[235]  =  14'b11000000100010;     //235pi/512
   cos[235]  =  14'b00001000001110;     //235pi/512
   sin[236]  =  14'b11000000011111;     //236pi/512
   cos[236]  =  14'b00000111110101;     //236pi/512
   sin[237]  =  14'b11000000011100;     //237pi/512
   cos[237]  =  14'b00000111011100;     //237pi/512
   sin[238]  =  14'b11000000011001;     //238pi/512
   cos[238]  =  14'b00000111000011;     //238pi/512
   sin[239]  =  14'b11000000010110;     //239pi/512
   cos[239]  =  14'b00000110101010;     //239pi/512
   sin[240]  =  14'b11000000010100;     //240pi/512
   cos[240]  =  14'b00000110010001;     //240pi/512
   sin[241]  =  14'b11000000010001;     //241pi/512
   cos[241]  =  14'b00000101111000;     //241pi/512
   sin[242]  =  14'b11000000001111;     //242pi/512
   cos[242]  =  14'b00000101011111;     //242pi/512
   sin[243]  =  14'b11000000001101;     //243pi/512
   cos[243]  =  14'b00000101000110;     //243pi/512
   sin[244]  =  14'b11000000001011;     //244pi/512
   cos[244]  =  14'b00000100101101;     //244pi/512
   sin[245]  =  14'b11000000001001;     //245pi/512
   cos[245]  =  14'b00000100010100;     //245pi/512
   sin[246]  =  14'b11000000001000;     //246pi/512
   cos[246]  =  14'b00000011111011;     //246pi/512
   sin[247]  =  14'b11000000000110;     //247pi/512
   cos[247]  =  14'b00000011100010;     //247pi/512
   sin[248]  =  14'b11000000000101;     //248pi/512
   cos[248]  =  14'b00000011001000;     //248pi/512
   sin[249]  =  14'b11000000000100;     //249pi/512
   cos[249]  =  14'b00000010101111;     //249pi/512
   sin[250]  =  14'b11000000000011;     //250pi/512
   cos[250]  =  14'b00000010010110;     //250pi/512
   sin[251]  =  14'b11000000000010;     //251pi/512
   cos[251]  =  14'b00000001111101;     //251pi/512
   sin[252]  =  14'b11000000000001;     //252pi/512
   cos[252]  =  14'b00000001100100;     //252pi/512
   sin[253]  =  14'b11000000000001;     //253pi/512
   cos[253]  =  14'b00000001001011;     //253pi/512
   sin[254]  =  14'b11000000000000;     //254pi/512
   cos[254]  =  14'b00000000110010;     //254pi/512
   sin[255]  =  14'b11000000000000;     //255pi/512
   cos[255]  =  14'b00000000011001;     //255pi/512
   sin[256]  =  14'b11000000000000;     //256pi/512
   cos[256]  =  14'b00000000000000;     //256pi/512
   sin[257]  =  14'b11000000000000;     //257pi/512
   cos[257]  =  14'b11111111100111;     //257pi/512
   sin[258]  =  14'b11000000000000;     //258pi/512
   cos[258]  =  14'b11111111001110;     //258pi/512
   sin[259]  =  14'b11000000000001;     //259pi/512
   cos[259]  =  14'b11111110110101;     //259pi/512
   sin[260]  =  14'b11000000000001;     //260pi/512
   cos[260]  =  14'b11111110011011;     //260pi/512
   sin[261]  =  14'b11000000000010;     //261pi/512
   cos[261]  =  14'b11111110000010;     //261pi/512
   sin[262]  =  14'b11000000000011;     //262pi/512
   cos[262]  =  14'b11111101101001;     //262pi/512
   sin[263]  =  14'b11000000000100;     //263pi/512
   cos[263]  =  14'b11111101010000;     //263pi/512
   sin[264]  =  14'b11000000000101;     //264pi/512
   cos[264]  =  14'b11111100110111;     //264pi/512
   sin[265]  =  14'b11000000000110;     //265pi/512
   cos[265]  =  14'b11111100011110;     //265pi/512
   sin[266]  =  14'b11000000001000;     //266pi/512
   cos[266]  =  14'b11111100000101;     //266pi/512
   sin[267]  =  14'b11000000001001;     //267pi/512
   cos[267]  =  14'b11111011101100;     //267pi/512
   sin[268]  =  14'b11000000001011;     //268pi/512
   cos[268]  =  14'b11111011010011;     //268pi/512
   sin[269]  =  14'b11000000001101;     //269pi/512
   cos[269]  =  14'b11111010111010;     //269pi/512
   sin[270]  =  14'b11000000001111;     //270pi/512
   cos[270]  =  14'b11111010100001;     //270pi/512
   sin[271]  =  14'b11000000010001;     //271pi/512
   cos[271]  =  14'b11111010001000;     //271pi/512
   sin[272]  =  14'b11000000010100;     //272pi/512
   cos[272]  =  14'b11111001101111;     //272pi/512
   sin[273]  =  14'b11000000010110;     //273pi/512
   cos[273]  =  14'b11111001010110;     //273pi/512
   sin[274]  =  14'b11000000011001;     //274pi/512
   cos[274]  =  14'b11111000111101;     //274pi/512
   sin[275]  =  14'b11000000011100;     //275pi/512
   cos[275]  =  14'b11111000100100;     //275pi/512
   sin[276]  =  14'b11000000011111;     //276pi/512
   cos[276]  =  14'b11111000001011;     //276pi/512
   sin[277]  =  14'b11000000100010;     //277pi/512
   cos[277]  =  14'b11110111110010;     //277pi/512
   sin[278]  =  14'b11000000100101;     //278pi/512
   cos[278]  =  14'b11110111011001;     //278pi/512
   sin[279]  =  14'b11000000101001;     //279pi/512
   cos[279]  =  14'b11110111000000;     //279pi/512
   sin[280]  =  14'b11000000101100;     //280pi/512
   cos[280]  =  14'b11110110100111;     //280pi/512
   sin[281]  =  14'b11000000110000;     //281pi/512
   cos[281]  =  14'b11110110001110;     //281pi/512
   sin[282]  =  14'b11000000110100;     //282pi/512
   cos[282]  =  14'b11110101110101;     //282pi/512
   sin[283]  =  14'b11000000111000;     //283pi/512
   cos[283]  =  14'b11110101011101;     //283pi/512
   sin[284]  =  14'b11000000111100;     //284pi/512
   cos[284]  =  14'b11110101000100;     //284pi/512
   sin[285]  =  14'b11000001000001;     //285pi/512
   cos[285]  =  14'b11110100101011;     //285pi/512
   sin[286]  =  14'b11000001000101;     //286pi/512
   cos[286]  =  14'b11110100010010;     //286pi/512
   sin[287]  =  14'b11000001001010;     //287pi/512
   cos[287]  =  14'b11110011111010;     //287pi/512
   sin[288]  =  14'b11000001001111;     //288pi/512
   cos[288]  =  14'b11110011100001;     //288pi/512
   sin[289]  =  14'b11000001010100;     //289pi/512
   cos[289]  =  14'b11110011001000;     //289pi/512
   sin[290]  =  14'b11000001011001;     //290pi/512
   cos[290]  =  14'b11110010110000;     //290pi/512
   sin[291]  =  14'b11000001011110;     //291pi/512
   cos[291]  =  14'b11110010010111;     //291pi/512
   sin[292]  =  14'b11000001100100;     //292pi/512
   cos[292]  =  14'b11110001111111;     //292pi/512
   sin[293]  =  14'b11000001101001;     //293pi/512
   cos[293]  =  14'b11110001100110;     //293pi/512
   sin[294]  =  14'b11000001101111;     //294pi/512
   cos[294]  =  14'b11110001001110;     //294pi/512
   sin[295]  =  14'b11000001110101;     //295pi/512
   cos[295]  =  14'b11110000110101;     //295pi/512
   sin[296]  =  14'b11000001111011;     //296pi/512
   cos[296]  =  14'b11110000011101;     //296pi/512
   sin[297]  =  14'b11000010000001;     //297pi/512
   cos[297]  =  14'b11110000000100;     //297pi/512
   sin[298]  =  14'b11000010000111;     //298pi/512
   cos[298]  =  14'b11101111101100;     //298pi/512
   sin[299]  =  14'b11000010001110;     //299pi/512
   cos[299]  =  14'b11101111010100;     //299pi/512
   sin[300]  =  14'b11000010010100;     //300pi/512
   cos[300]  =  14'b11101110111100;     //300pi/512
   sin[301]  =  14'b11000010011011;     //301pi/512
   cos[301]  =  14'b11101110100011;     //301pi/512
   sin[302]  =  14'b11000010100010;     //302pi/512
   cos[302]  =  14'b11101110001011;     //302pi/512
   sin[303]  =  14'b11000010101001;     //303pi/512
   cos[303]  =  14'b11101101110011;     //303pi/512
   sin[304]  =  14'b11000010110000;     //304pi/512
   cos[304]  =  14'b11101101011011;     //304pi/512
   sin[305]  =  14'b11000010111000;     //305pi/512
   cos[305]  =  14'b11101101000011;     //305pi/512
   sin[306]  =  14'b11000010111111;     //306pi/512
   cos[306]  =  14'b11101100101011;     //306pi/512
   sin[307]  =  14'b11000011000111;     //307pi/512
   cos[307]  =  14'b11101100010011;     //307pi/512
   sin[308]  =  14'b11000011001111;     //308pi/512
   cos[308]  =  14'b11101011111011;     //308pi/512
   sin[309]  =  14'b11000011010111;     //309pi/512
   cos[309]  =  14'b11101011100011;     //309pi/512
   sin[310]  =  14'b11000011011111;     //310pi/512
   cos[310]  =  14'b11101011001100;     //310pi/512
   sin[311]  =  14'b11000011100111;     //311pi/512
   cos[311]  =  14'b11101010110100;     //311pi/512
   sin[312]  =  14'b11000011101111;     //312pi/512
   cos[312]  =  14'b11101010011100;     //312pi/512
   sin[313]  =  14'b11000011111000;     //313pi/512
   cos[313]  =  14'b11101010000100;     //313pi/512
   sin[314]  =  14'b11000100000001;     //314pi/512
   cos[314]  =  14'b11101001101101;     //314pi/512
   sin[315]  =  14'b11000100001001;     //315pi/512
   cos[315]  =  14'b11101001010101;     //315pi/512
   sin[316]  =  14'b11000100010010;     //316pi/512
   cos[316]  =  14'b11101000111110;     //316pi/512
   sin[317]  =  14'b11000100011100;     //317pi/512
   cos[317]  =  14'b11101000100110;     //317pi/512
   sin[318]  =  14'b11000100100101;     //318pi/512
   cos[318]  =  14'b11101000001111;     //318pi/512
   sin[319]  =  14'b11000100101110;     //319pi/512
   cos[319]  =  14'b11100111111000;     //319pi/512
   sin[320]  =  14'b11000100111000;     //320pi/512
   cos[320]  =  14'b11100111100001;     //320pi/512
   sin[321]  =  14'b11000101000001;     //321pi/512
   cos[321]  =  14'b11100111001001;     //321pi/512
   sin[322]  =  14'b11000101001011;     //322pi/512
   cos[322]  =  14'b11100110110010;     //322pi/512
   sin[323]  =  14'b11000101010101;     //323pi/512
   cos[323]  =  14'b11100110011011;     //323pi/512
   sin[324]  =  14'b11000101011111;     //324pi/512
   cos[324]  =  14'b11100110000100;     //324pi/512
   sin[325]  =  14'b11000101101010;     //325pi/512
   cos[325]  =  14'b11100101101101;     //325pi/512
   sin[326]  =  14'b11000101110100;     //326pi/512
   cos[326]  =  14'b11100101010110;     //326pi/512
   sin[327]  =  14'b11000101111111;     //327pi/512
   cos[327]  =  14'b11100100111111;     //327pi/512
   sin[328]  =  14'b11000110001001;     //328pi/512
   cos[328]  =  14'b11100100101001;     //328pi/512
   sin[329]  =  14'b11000110010100;     //329pi/512
   cos[329]  =  14'b11100100010010;     //329pi/512
   sin[330]  =  14'b11000110011111;     //330pi/512
   cos[330]  =  14'b11100011111011;     //330pi/512
   sin[331]  =  14'b11000110101010;     //331pi/512
   cos[331]  =  14'b11100011100101;     //331pi/512
   sin[332]  =  14'b11000110110101;     //332pi/512
   cos[332]  =  14'b11100011001110;     //332pi/512
   sin[333]  =  14'b11000111000001;     //333pi/512
   cos[333]  =  14'b11100010111000;     //333pi/512
   sin[334]  =  14'b11000111001100;     //334pi/512
   cos[334]  =  14'b11100010100010;     //334pi/512
   sin[335]  =  14'b11000111011000;     //335pi/512
   cos[335]  =  14'b11100010001011;     //335pi/512
   sin[336]  =  14'b11000111100100;     //336pi/512
   cos[336]  =  14'b11100001110101;     //336pi/512
   sin[337]  =  14'b11000111110000;     //337pi/512
   cos[337]  =  14'b11100001011111;     //337pi/512
   sin[338]  =  14'b11000111111100;     //338pi/512
   cos[338]  =  14'b11100001001001;     //338pi/512
   sin[339]  =  14'b11001000001000;     //339pi/512
   cos[339]  =  14'b11100000110011;     //339pi/512
   sin[340]  =  14'b11001000010100;     //340pi/512
   cos[340]  =  14'b11100000011101;     //340pi/512
   sin[341]  =  14'b11001000100001;     //341pi/512
   cos[341]  =  14'b11100000000111;     //341pi/512
   sin[342]  =  14'b11001000101101;     //342pi/512
   cos[342]  =  14'b11011111110010;     //342pi/512
   sin[343]  =  14'b11001000111010;     //343pi/512
   cos[343]  =  14'b11011111011100;     //343pi/512
   sin[344]  =  14'b11001001000111;     //344pi/512
   cos[344]  =  14'b11011111000110;     //344pi/512
   sin[345]  =  14'b11001001010100;     //345pi/512
   cos[345]  =  14'b11011110110001;     //345pi/512
   sin[346]  =  14'b11001001100001;     //346pi/512
   cos[346]  =  14'b11011110011011;     //346pi/512
   sin[347]  =  14'b11001001101110;     //347pi/512
   cos[347]  =  14'b11011110000110;     //347pi/512
   sin[348]  =  14'b11001001111011;     //348pi/512
   cos[348]  =  14'b11011101110001;     //348pi/512
   sin[349]  =  14'b11001010001001;     //349pi/512
   cos[349]  =  14'b11011101011011;     //349pi/512
   sin[350]  =  14'b11001010010111;     //350pi/512
   cos[350]  =  14'b11011101000110;     //350pi/512
   sin[351]  =  14'b11001010100100;     //351pi/512
   cos[351]  =  14'b11011100110001;     //351pi/512
   sin[352]  =  14'b11001010110010;     //352pi/512
   cos[352]  =  14'b11011100011100;     //352pi/512
   sin[353]  =  14'b11001011000000;     //353pi/512
   cos[353]  =  14'b11011100001000;     //353pi/512
   sin[354]  =  14'b11001011001110;     //354pi/512
   cos[354]  =  14'b11011011110011;     //354pi/512
   sin[355]  =  14'b11001011011101;     //355pi/512
   cos[355]  =  14'b11011011011110;     //355pi/512
   sin[356]  =  14'b11001011101011;     //356pi/512
   cos[356]  =  14'b11011011001001;     //356pi/512
   sin[357]  =  14'b11001011111010;     //357pi/512
   cos[357]  =  14'b11011010110101;     //357pi/512
   sin[358]  =  14'b11001100001000;     //358pi/512
   cos[358]  =  14'b11011010100001;     //358pi/512
   sin[359]  =  14'b11001100010111;     //359pi/512
   cos[359]  =  14'b11011010001100;     //359pi/512
   sin[360]  =  14'b11001100100110;     //360pi/512
   cos[360]  =  14'b11011001111000;     //360pi/512
   sin[361]  =  14'b11001100110101;     //361pi/512
   cos[361]  =  14'b11011001100100;     //361pi/512
   sin[362]  =  14'b11001101000100;     //362pi/512
   cos[362]  =  14'b11011001010000;     //362pi/512
   sin[363]  =  14'b11001101010100;     //363pi/512
   cos[363]  =  14'b11011000111100;     //363pi/512
   sin[364]  =  14'b11001101100011;     //364pi/512
   cos[364]  =  14'b11011000101000;     //364pi/512
   sin[365]  =  14'b11001101110010;     //365pi/512
   cos[365]  =  14'b11011000010100;     //365pi/512
   sin[366]  =  14'b11001110000010;     //366pi/512
   cos[366]  =  14'b11011000000001;     //366pi/512
   sin[367]  =  14'b11001110010010;     //367pi/512
   cos[367]  =  14'b11010111101101;     //367pi/512
   sin[368]  =  14'b11001110100010;     //368pi/512
   cos[368]  =  14'b11010111011010;     //368pi/512
   sin[369]  =  14'b11001110110010;     //369pi/512
   cos[369]  =  14'b11010111000110;     //369pi/512
   sin[370]  =  14'b11001111000010;     //370pi/512
   cos[370]  =  14'b11010110110011;     //370pi/512
   sin[371]  =  14'b11001111010010;     //371pi/512
   cos[371]  =  14'b11010110100000;     //371pi/512
   sin[372]  =  14'b11001111100010;     //372pi/512
   cos[372]  =  14'b11010110001101;     //372pi/512
   sin[373]  =  14'b11001111110011;     //373pi/512
   cos[373]  =  14'b11010101111010;     //373pi/512
   sin[374]  =  14'b11010000000100;     //374pi/512
   cos[374]  =  14'b11010101100111;     //374pi/512
   sin[375]  =  14'b11010000010100;     //375pi/512
   cos[375]  =  14'b11010101010100;     //375pi/512
   sin[376]  =  14'b11010000100101;     //376pi/512
   cos[376]  =  14'b11010101000001;     //376pi/512
   sin[377]  =  14'b11010000110110;     //377pi/512
   cos[377]  =  14'b11010100101111;     //377pi/512
   sin[378]  =  14'b11010001000111;     //378pi/512
   cos[378]  =  14'b11010100011100;     //378pi/512
   sin[379]  =  14'b11010001011000;     //379pi/512
   cos[379]  =  14'b11010100001010;     //379pi/512
   sin[380]  =  14'b11010001101001;     //380pi/512
   cos[380]  =  14'b11010011111000;     //380pi/512
   sin[381]  =  14'b11010001111011;     //381pi/512
   cos[381]  =  14'b11010011100101;     //381pi/512
   sin[382]  =  14'b11010010001100;     //382pi/512
   cos[382]  =  14'b11010011010011;     //382pi/512
   sin[383]  =  14'b11010010011110;     //383pi/512
   cos[383]  =  14'b11010011000010;     //383pi/512
   sin[384]  =  14'b11010010110000;     //384pi/512
   cos[384]  =  14'b11010010110000;     //384pi/512
   sin[385]  =  14'b11010011000010;     //385pi/512
   cos[385]  =  14'b11010010011110;     //385pi/512
   sin[386]  =  14'b11010011010011;     //386pi/512
   cos[386]  =  14'b11010010001100;     //386pi/512
   sin[387]  =  14'b11010011100101;     //387pi/512
   cos[387]  =  14'b11010001111011;     //387pi/512
   sin[388]  =  14'b11010011111000;     //388pi/512
   cos[388]  =  14'b11010001101001;     //388pi/512
   sin[389]  =  14'b11010100001010;     //389pi/512
   cos[389]  =  14'b11010001011000;     //389pi/512
   sin[390]  =  14'b11010100011100;     //390pi/512
   cos[390]  =  14'b11010001000111;     //390pi/512
   sin[391]  =  14'b11010100101111;     //391pi/512
   cos[391]  =  14'b11010000110110;     //391pi/512
   sin[392]  =  14'b11010101000001;     //392pi/512
   cos[392]  =  14'b11010000100101;     //392pi/512
   sin[393]  =  14'b11010101010100;     //393pi/512
   cos[393]  =  14'b11010000010100;     //393pi/512
   sin[394]  =  14'b11010101100111;     //394pi/512
   cos[394]  =  14'b11010000000100;     //394pi/512
   sin[395]  =  14'b11010101111010;     //395pi/512
   cos[395]  =  14'b11001111110011;     //395pi/512
   sin[396]  =  14'b11010110001101;     //396pi/512
   cos[396]  =  14'b11001111100010;     //396pi/512
   sin[397]  =  14'b11010110100000;     //397pi/512
   cos[397]  =  14'b11001111010010;     //397pi/512
   sin[398]  =  14'b11010110110011;     //398pi/512
   cos[398]  =  14'b11001111000010;     //398pi/512
   sin[399]  =  14'b11010111000110;     //399pi/512
   cos[399]  =  14'b11001110110010;     //399pi/512
   sin[400]  =  14'b11010111011010;     //400pi/512
   cos[400]  =  14'b11001110100010;     //400pi/512
   sin[401]  =  14'b11010111101101;     //401pi/512
   cos[401]  =  14'b11001110010010;     //401pi/512
   sin[402]  =  14'b11011000000001;     //402pi/512
   cos[402]  =  14'b11001110000010;     //402pi/512
   sin[403]  =  14'b11011000010100;     //403pi/512
   cos[403]  =  14'b11001101110010;     //403pi/512
   sin[404]  =  14'b11011000101000;     //404pi/512
   cos[404]  =  14'b11001101100011;     //404pi/512
   sin[405]  =  14'b11011000111100;     //405pi/512
   cos[405]  =  14'b11001101010100;     //405pi/512
   sin[406]  =  14'b11011001010000;     //406pi/512
   cos[406]  =  14'b11001101000100;     //406pi/512
   sin[407]  =  14'b11011001100100;     //407pi/512
   cos[407]  =  14'b11001100110101;     //407pi/512
   sin[408]  =  14'b11011001111000;     //408pi/512
   cos[408]  =  14'b11001100100110;     //408pi/512
   sin[409]  =  14'b11011010001100;     //409pi/512
   cos[409]  =  14'b11001100010111;     //409pi/512
   sin[410]  =  14'b11011010100001;     //410pi/512
   cos[410]  =  14'b11001100001000;     //410pi/512
   sin[411]  =  14'b11011010110101;     //411pi/512
   cos[411]  =  14'b11001011111010;     //411pi/512
   sin[412]  =  14'b11011011001001;     //412pi/512
   cos[412]  =  14'b11001011101011;     //412pi/512
   sin[413]  =  14'b11011011011110;     //413pi/512
   cos[413]  =  14'b11001011011101;     //413pi/512
   sin[414]  =  14'b11011011110011;     //414pi/512
   cos[414]  =  14'b11001011001110;     //414pi/512
   sin[415]  =  14'b11011100001000;     //415pi/512
   cos[415]  =  14'b11001011000000;     //415pi/512
   sin[416]  =  14'b11011100011100;     //416pi/512
   cos[416]  =  14'b11001010110010;     //416pi/512
   sin[417]  =  14'b11011100110001;     //417pi/512
   cos[417]  =  14'b11001010100100;     //417pi/512
   sin[418]  =  14'b11011101000110;     //418pi/512
   cos[418]  =  14'b11001010010111;     //418pi/512
   sin[419]  =  14'b11011101011011;     //419pi/512
   cos[419]  =  14'b11001010001001;     //419pi/512
   sin[420]  =  14'b11011101110001;     //420pi/512
   cos[420]  =  14'b11001001111011;     //420pi/512
   sin[421]  =  14'b11011110000110;     //421pi/512
   cos[421]  =  14'b11001001101110;     //421pi/512
   sin[422]  =  14'b11011110011011;     //422pi/512
   cos[422]  =  14'b11001001100001;     //422pi/512
   sin[423]  =  14'b11011110110001;     //423pi/512
   cos[423]  =  14'b11001001010100;     //423pi/512
   sin[424]  =  14'b11011111000110;     //424pi/512
   cos[424]  =  14'b11001001000111;     //424pi/512
   sin[425]  =  14'b11011111011100;     //425pi/512
   cos[425]  =  14'b11001000111010;     //425pi/512
   sin[426]  =  14'b11011111110010;     //426pi/512
   cos[426]  =  14'b11001000101101;     //426pi/512
   sin[427]  =  14'b11100000000111;     //427pi/512
   cos[427]  =  14'b11001000100001;     //427pi/512
   sin[428]  =  14'b11100000011101;     //428pi/512
   cos[428]  =  14'b11001000010100;     //428pi/512
   sin[429]  =  14'b11100000110011;     //429pi/512
   cos[429]  =  14'b11001000001000;     //429pi/512
   sin[430]  =  14'b11100001001001;     //430pi/512
   cos[430]  =  14'b11000111111100;     //430pi/512
   sin[431]  =  14'b11100001011111;     //431pi/512
   cos[431]  =  14'b11000111110000;     //431pi/512
   sin[432]  =  14'b11100001110101;     //432pi/512
   cos[432]  =  14'b11000111100100;     //432pi/512
   sin[433]  =  14'b11100010001011;     //433pi/512
   cos[433]  =  14'b11000111011000;     //433pi/512
   sin[434]  =  14'b11100010100010;     //434pi/512
   cos[434]  =  14'b11000111001100;     //434pi/512
   sin[435]  =  14'b11100010111000;     //435pi/512
   cos[435]  =  14'b11000111000001;     //435pi/512
   sin[436]  =  14'b11100011001110;     //436pi/512
   cos[436]  =  14'b11000110110101;     //436pi/512
   sin[437]  =  14'b11100011100101;     //437pi/512
   cos[437]  =  14'b11000110101010;     //437pi/512
   sin[438]  =  14'b11100011111011;     //438pi/512
   cos[438]  =  14'b11000110011111;     //438pi/512
   sin[439]  =  14'b11100100010010;     //439pi/512
   cos[439]  =  14'b11000110010100;     //439pi/512
   sin[440]  =  14'b11100100101001;     //440pi/512
   cos[440]  =  14'b11000110001001;     //440pi/512
   sin[441]  =  14'b11100100111111;     //441pi/512
   cos[441]  =  14'b11000101111111;     //441pi/512
   sin[442]  =  14'b11100101010110;     //442pi/512
   cos[442]  =  14'b11000101110100;     //442pi/512
   sin[443]  =  14'b11100101101101;     //443pi/512
   cos[443]  =  14'b11000101101010;     //443pi/512
   sin[444]  =  14'b11100110000100;     //444pi/512
   cos[444]  =  14'b11000101011111;     //444pi/512
   sin[445]  =  14'b11100110011011;     //445pi/512
   cos[445]  =  14'b11000101010101;     //445pi/512
   sin[446]  =  14'b11100110110010;     //446pi/512
   cos[446]  =  14'b11000101001011;     //446pi/512
   sin[447]  =  14'b11100111001001;     //447pi/512
   cos[447]  =  14'b11000101000001;     //447pi/512
   sin[448]  =  14'b11100111100001;     //448pi/512
   cos[448]  =  14'b11000100111000;     //448pi/512
   sin[449]  =  14'b11100111111000;     //449pi/512
   cos[449]  =  14'b11000100101110;     //449pi/512
   sin[450]  =  14'b11101000001111;     //450pi/512
   cos[450]  =  14'b11000100100101;     //450pi/512
   sin[451]  =  14'b11101000100110;     //451pi/512
   cos[451]  =  14'b11000100011100;     //451pi/512
   sin[452]  =  14'b11101000111110;     //452pi/512
   cos[452]  =  14'b11000100010010;     //452pi/512
   sin[453]  =  14'b11101001010101;     //453pi/512
   cos[453]  =  14'b11000100001001;     //453pi/512
   sin[454]  =  14'b11101001101101;     //454pi/512
   cos[454]  =  14'b11000100000001;     //454pi/512
   sin[455]  =  14'b11101010000100;     //455pi/512
   cos[455]  =  14'b11000011111000;     //455pi/512
   sin[456]  =  14'b11101010011100;     //456pi/512
   cos[456]  =  14'b11000011101111;     //456pi/512
   sin[457]  =  14'b11101010110100;     //457pi/512
   cos[457]  =  14'b11000011100111;     //457pi/512
   sin[458]  =  14'b11101011001100;     //458pi/512
   cos[458]  =  14'b11000011011111;     //458pi/512
   sin[459]  =  14'b11101011100011;     //459pi/512
   cos[459]  =  14'b11000011010111;     //459pi/512
   sin[460]  =  14'b11101011111011;     //460pi/512
   cos[460]  =  14'b11000011001111;     //460pi/512
   sin[461]  =  14'b11101100010011;     //461pi/512
   cos[461]  =  14'b11000011000111;     //461pi/512
   sin[462]  =  14'b11101100101011;     //462pi/512
   cos[462]  =  14'b11000010111111;     //462pi/512
   sin[463]  =  14'b11101101000011;     //463pi/512
   cos[463]  =  14'b11000010111000;     //463pi/512
   sin[464]  =  14'b11101101011011;     //464pi/512
   cos[464]  =  14'b11000010110000;     //464pi/512
   sin[465]  =  14'b11101101110011;     //465pi/512
   cos[465]  =  14'b11000010101001;     //465pi/512
   sin[466]  =  14'b11101110001011;     //466pi/512
   cos[466]  =  14'b11000010100010;     //466pi/512
   sin[467]  =  14'b11101110100011;     //467pi/512
   cos[467]  =  14'b11000010011011;     //467pi/512
   sin[468]  =  14'b11101110111100;     //468pi/512
   cos[468]  =  14'b11000010010100;     //468pi/512
   sin[469]  =  14'b11101111010100;     //469pi/512
   cos[469]  =  14'b11000010001110;     //469pi/512
   sin[470]  =  14'b11101111101100;     //470pi/512
   cos[470]  =  14'b11000010000111;     //470pi/512
   sin[471]  =  14'b11110000000100;     //471pi/512
   cos[471]  =  14'b11000010000001;     //471pi/512
   sin[472]  =  14'b11110000011101;     //472pi/512
   cos[472]  =  14'b11000001111011;     //472pi/512
   sin[473]  =  14'b11110000110101;     //473pi/512
   cos[473]  =  14'b11000001110101;     //473pi/512
   sin[474]  =  14'b11110001001110;     //474pi/512
   cos[474]  =  14'b11000001101111;     //474pi/512
   sin[475]  =  14'b11110001100110;     //475pi/512
   cos[475]  =  14'b11000001101001;     //475pi/512
   sin[476]  =  14'b11110001111111;     //476pi/512
   cos[476]  =  14'b11000001100100;     //476pi/512
   sin[477]  =  14'b11110010010111;     //477pi/512
   cos[477]  =  14'b11000001011110;     //477pi/512
   sin[478]  =  14'b11110010110000;     //478pi/512
   cos[478]  =  14'b11000001011001;     //478pi/512
   sin[479]  =  14'b11110011001000;     //479pi/512
   cos[479]  =  14'b11000001010100;     //479pi/512
   sin[480]  =  14'b11110011100001;     //480pi/512
   cos[480]  =  14'b11000001001111;     //480pi/512
   sin[481]  =  14'b11110011111010;     //481pi/512
   cos[481]  =  14'b11000001001010;     //481pi/512
   sin[482]  =  14'b11110100010010;     //482pi/512
   cos[482]  =  14'b11000001000101;     //482pi/512
   sin[483]  =  14'b11110100101011;     //483pi/512
   cos[483]  =  14'b11000001000001;     //483pi/512
   sin[484]  =  14'b11110101000100;     //484pi/512
   cos[484]  =  14'b11000000111100;     //484pi/512
   sin[485]  =  14'b11110101011101;     //485pi/512
   cos[485]  =  14'b11000000111000;     //485pi/512
   sin[486]  =  14'b11110101110101;     //486pi/512
   cos[486]  =  14'b11000000110100;     //486pi/512
   sin[487]  =  14'b11110110001110;     //487pi/512
   cos[487]  =  14'b11000000110000;     //487pi/512
   sin[488]  =  14'b11110110100111;     //488pi/512
   cos[488]  =  14'b11000000101100;     //488pi/512
   sin[489]  =  14'b11110111000000;     //489pi/512
   cos[489]  =  14'b11000000101001;     //489pi/512
   sin[490]  =  14'b11110111011001;     //490pi/512
   cos[490]  =  14'b11000000100101;     //490pi/512
   sin[491]  =  14'b11110111110010;     //491pi/512
   cos[491]  =  14'b11000000100010;     //491pi/512
   sin[492]  =  14'b11111000001011;     //492pi/512
   cos[492]  =  14'b11000000011111;     //492pi/512
   sin[493]  =  14'b11111000100100;     //493pi/512
   cos[493]  =  14'b11000000011100;     //493pi/512
   sin[494]  =  14'b11111000111101;     //494pi/512
   cos[494]  =  14'b11000000011001;     //494pi/512
   sin[495]  =  14'b11111001010110;     //495pi/512
   cos[495]  =  14'b11000000010110;     //495pi/512
   sin[496]  =  14'b11111001101111;     //496pi/512
   cos[496]  =  14'b11000000010100;     //496pi/512
   sin[497]  =  14'b11111010001000;     //497pi/512
   cos[497]  =  14'b11000000010001;     //497pi/512
   sin[498]  =  14'b11111010100001;     //498pi/512
   cos[498]  =  14'b11000000001111;     //498pi/512
   sin[499]  =  14'b11111010111010;     //499pi/512
   cos[499]  =  14'b11000000001101;     //499pi/512
   sin[500]  =  14'b11111011010011;     //500pi/512
   cos[500]  =  14'b11000000001011;     //500pi/512
   sin[501]  =  14'b11111011101100;     //501pi/512
   cos[501]  =  14'b11000000001001;     //501pi/512
   sin[502]  =  14'b11111100000101;     //502pi/512
   cos[502]  =  14'b11000000001000;     //502pi/512
   sin[503]  =  14'b11111100011110;     //503pi/512
   cos[503]  =  14'b11000000000110;     //503pi/512
   sin[504]  =  14'b11111100110111;     //504pi/512
   cos[504]  =  14'b11000000000101;     //504pi/512
   sin[505]  =  14'b11111101010000;     //505pi/512
   cos[505]  =  14'b11000000000100;     //505pi/512
   sin[506]  =  14'b11111101101001;     //506pi/512
   cos[506]  =  14'b11000000000011;     //506pi/512
   sin[507]  =  14'b11111110000010;     //507pi/512
   cos[507]  =  14'b11000000000010;     //507pi/512
   sin[508]  =  14'b11111110011011;     //508pi/512
   cos[508]  =  14'b11000000000001;     //508pi/512
   sin[509]  =  14'b11111110110101;     //509pi/512
   cos[509]  =  14'b11000000000001;     //509pi/512
   sin[510]  =  14'b11111111001110;     //510pi/512
   cos[510]  =  14'b11000000000000;     //510pi/512
   sin[511]  =  14'b11111111100111;     //511pi/512
   cos[511]  =  14'b11000000000000;     //511pi/512

///////////////////////////////////////////////////////////////
   m_sin[0]  =  14'b00000000000000;     //0pi/512
   m_cos[0]  =  14'b01000000000000;     //0pi/512
   m_sin[1]  =  14'b11111111101011;     //1pi/512
   m_cos[1]  =  14'b00111111111111;     //1pi/512
   m_sin[2]  =  14'b11111111010101;     //2pi/512
   m_cos[2]  =  14'b00111111111111;     //2pi/512
   m_sin[3]  =  14'b11111111000000;     //3pi/512
   m_cos[3]  =  14'b00111111111111;     //3pi/512
   m_sin[4]  =  14'b11111110101011;     //4pi/512
   m_cos[4]  =  14'b00111111111111;     //4pi/512
   m_sin[5]  =  14'b11111110010101;     //5pi/512
   m_cos[5]  =  14'b00111111111110;     //5pi/512
   m_sin[6]  =  14'b11111110000000;     //6pi/512
   m_cos[6]  =  14'b00111111111101;     //6pi/512
   m_sin[7]  =  14'b11111101101010;     //7pi/512
   m_cos[7]  =  14'b00111111111101;     //7pi/512
   m_sin[8]  =  14'b11111101010101;     //8pi/512
   m_cos[8]  =  14'b00111111111100;     //8pi/512
   m_sin[9]  =  14'b11111101000000;     //9pi/512
   m_cos[9]  =  14'b00111111111011;     //9pi/512
   m_sin[10]  =  14'b11111100101010;     //10pi/512
   m_cos[10]  =  14'b00111111111010;     //10pi/512
   m_sin[11]  =  14'b11111100010101;     //11pi/512
   m_cos[11]  =  14'b00111111111001;     //11pi/512
   m_sin[12]  =  14'b11111100000000;     //12pi/512
   m_cos[12]  =  14'b00111111110111;     //12pi/512
   m_sin[13]  =  14'b11111011101010;     //13pi/512
   m_cos[13]  =  14'b00111111110110;     //13pi/512
   m_sin[14]  =  14'b11111011010101;     //14pi/512
   m_cos[14]  =  14'b00111111110101;     //14pi/512
   m_sin[15]  =  14'b11111011000000;     //15pi/512
   m_cos[15]  =  14'b00111111110011;     //15pi/512
   m_sin[16]  =  14'b11111010101011;     //16pi/512
   m_cos[16]  =  14'b00111111110001;     //16pi/512
   m_sin[17]  =  14'b11111010010101;     //17pi/512
   m_cos[17]  =  14'b00111111101111;     //17pi/512
   m_sin[18]  =  14'b11111010000000;     //18pi/512
   m_cos[18]  =  14'b00111111101101;     //18pi/512
   m_sin[19]  =  14'b11111001101011;     //19pi/512
   m_cos[19]  =  14'b00111111101011;     //19pi/512
   m_sin[20]  =  14'b11111001010110;     //20pi/512
   m_cos[20]  =  14'b00111111101001;     //20pi/512
   m_sin[21]  =  14'b11111001000000;     //21pi/512
   m_cos[21]  =  14'b00111111100111;     //21pi/512
   m_sin[22]  =  14'b11111000101011;     //22pi/512
   m_cos[22]  =  14'b00111111100101;     //22pi/512
   m_sin[23]  =  14'b11111000010110;     //23pi/512
   m_cos[23]  =  14'b00111111100010;     //23pi/512
   m_sin[24]  =  14'b11111000000001;     //24pi/512
   m_cos[24]  =  14'b00111111011111;     //24pi/512
   m_sin[25]  =  14'b11110111101011;     //25pi/512
   m_cos[25]  =  14'b00111111011101;     //25pi/512
   m_sin[26]  =  14'b11110111010110;     //26pi/512
   m_cos[26]  =  14'b00111111011010;     //26pi/512
   m_sin[27]  =  14'b11110111000001;     //27pi/512
   m_cos[27]  =  14'b00111111010111;     //27pi/512
   m_sin[28]  =  14'b11110110101100;     //28pi/512
   m_cos[28]  =  14'b00111111010100;     //28pi/512
   m_sin[29]  =  14'b11110110010111;     //29pi/512
   m_cos[29]  =  14'b00111111010001;     //29pi/512
   m_sin[30]  =  14'b11110110000010;     //30pi/512
   m_cos[30]  =  14'b00111111001101;     //30pi/512
   m_sin[31]  =  14'b11110101101101;     //31pi/512
   m_cos[31]  =  14'b00111111001010;     //31pi/512
   m_sin[32]  =  14'b11110101011000;     //32pi/512
   m_cos[32]  =  14'b00111111000111;     //32pi/512
   m_sin[33]  =  14'b11110101000011;     //33pi/512
   m_cos[33]  =  14'b00111111000011;     //33pi/512
   m_sin[34]  =  14'b11110100101101;     //34pi/512
   m_cos[34]  =  14'b00111110111111;     //34pi/512
   m_sin[35]  =  14'b11110100011000;     //35pi/512
   m_cos[35]  =  14'b00111110111011;     //35pi/512
   m_sin[36]  =  14'b11110100000011;     //36pi/512
   m_cos[36]  =  14'b00111110111000;     //36pi/512
   m_sin[37]  =  14'b11110011101110;     //37pi/512
   m_cos[37]  =  14'b00111110110011;     //37pi/512
   m_sin[38]  =  14'b11110011011010;     //38pi/512
   m_cos[38]  =  14'b00111110101111;     //38pi/512
   m_sin[39]  =  14'b11110011000101;     //39pi/512
   m_cos[39]  =  14'b00111110101011;     //39pi/512
   m_sin[40]  =  14'b11110010110000;     //40pi/512
   m_cos[40]  =  14'b00111110100111;     //40pi/512
   m_sin[41]  =  14'b11110010011011;     //41pi/512
   m_cos[41]  =  14'b00111110100010;     //41pi/512
   m_sin[42]  =  14'b11110010000110;     //42pi/512
   m_cos[42]  =  14'b00111110011110;     //42pi/512
   m_sin[43]  =  14'b11110001110001;     //43pi/512
   m_cos[43]  =  14'b00111110011001;     //43pi/512
   m_sin[44]  =  14'b11110001011100;     //44pi/512
   m_cos[44]  =  14'b00111110010100;     //44pi/512
   m_sin[45]  =  14'b11110001000111;     //45pi/512
   m_cos[45]  =  14'b00111110001111;     //45pi/512
   m_sin[46]  =  14'b11110000110011;     //46pi/512
   m_cos[46]  =  14'b00111110001010;     //46pi/512
   m_sin[47]  =  14'b11110000011110;     //47pi/512
   m_cos[47]  =  14'b00111110000101;     //47pi/512
   m_sin[48]  =  14'b11110000001001;     //48pi/512
   m_cos[48]  =  14'b00111110000000;     //48pi/512
   m_sin[49]  =  14'b11101111110101;     //49pi/512
   m_cos[49]  =  14'b00111101111010;     //49pi/512
   m_sin[50]  =  14'b11101111100000;     //50pi/512
   m_cos[50]  =  14'b00111101110101;     //50pi/512
   m_sin[51]  =  14'b11101111001011;     //51pi/512
   m_cos[51]  =  14'b00111101101111;     //51pi/512
   m_sin[52]  =  14'b11101110110111;     //52pi/512
   m_cos[52]  =  14'b00111101101010;     //52pi/512
   m_sin[53]  =  14'b11101110100010;     //53pi/512
   m_cos[53]  =  14'b00111101100100;     //53pi/512
   m_sin[54]  =  14'b11101110001110;     //54pi/512
   m_cos[54]  =  14'b00111101011110;     //54pi/512
   m_sin[55]  =  14'b11101101111001;     //55pi/512
   m_cos[55]  =  14'b00111101011000;     //55pi/512
   m_sin[56]  =  14'b11101101100101;     //56pi/512
   m_cos[56]  =  14'b00111101010010;     //56pi/512
   m_sin[57]  =  14'b11101101010000;     //57pi/512
   m_cos[57]  =  14'b00111101001100;     //57pi/512
   m_sin[58]  =  14'b11101100111100;     //58pi/512
   m_cos[58]  =  14'b00111101000110;     //58pi/512
   m_sin[59]  =  14'b11101100100111;     //59pi/512
   m_cos[59]  =  14'b00111100111111;     //59pi/512
   m_sin[60]  =  14'b11101100010011;     //60pi/512
   m_cos[60]  =  14'b00111100111001;     //60pi/512
   m_sin[61]  =  14'b11101011111111;     //61pi/512
   m_cos[61]  =  14'b00111100110010;     //61pi/512
   m_sin[62]  =  14'b11101011101010;     //62pi/512
   m_cos[62]  =  14'b00111100101011;     //62pi/512
   m_sin[63]  =  14'b11101011010110;     //63pi/512
   m_cos[63]  =  14'b00111100100100;     //63pi/512
   m_sin[64]  =  14'b11101011000010;     //64pi/512
   m_cos[64]  =  14'b00111100011101;     //64pi/512
   m_sin[65]  =  14'b11101010101110;     //65pi/512
   m_cos[65]  =  14'b00111100010110;     //65pi/512
   m_sin[66]  =  14'b11101010011010;     //66pi/512
   m_cos[66]  =  14'b00111100001111;     //66pi/512
   m_sin[67]  =  14'b11101010000110;     //67pi/512
   m_cos[67]  =  14'b00111100001000;     //67pi/512
   m_sin[68]  =  14'b11101001110010;     //68pi/512
   m_cos[68]  =  14'b00111100000001;     //68pi/512
   m_sin[69]  =  14'b11101001011110;     //69pi/512
   m_cos[69]  =  14'b00111011111001;     //69pi/512
   m_sin[70]  =  14'b11101001001010;     //70pi/512
   m_cos[70]  =  14'b00111011110010;     //70pi/512
   m_sin[71]  =  14'b11101000110110;     //71pi/512
   m_cos[71]  =  14'b00111011101010;     //71pi/512
   m_sin[72]  =  14'b11101000100010;     //72pi/512
   m_cos[72]  =  14'b00111011100010;     //72pi/512
   m_sin[73]  =  14'b11101000001110;     //73pi/512
   m_cos[73]  =  14'b00111011011010;     //73pi/512
   m_sin[74]  =  14'b11100111111010;     //74pi/512
   m_cos[74]  =  14'b00111011010010;     //74pi/512
   m_sin[75]  =  14'b11100111100110;     //75pi/512
   m_cos[75]  =  14'b00111011001010;     //75pi/512
   m_sin[76]  =  14'b11100111010011;     //76pi/512
   m_cos[76]  =  14'b00111011000010;     //76pi/512
   m_sin[77]  =  14'b11100110111111;     //77pi/512
   m_cos[77]  =  14'b00111010111010;     //77pi/512
   m_sin[78]  =  14'b11100110101011;     //78pi/512
   m_cos[78]  =  14'b00111010110001;     //78pi/512
   m_sin[79]  =  14'b11100110011000;     //79pi/512
   m_cos[79]  =  14'b00111010101001;     //79pi/512
   m_sin[80]  =  14'b11100110000100;     //80pi/512
   m_cos[80]  =  14'b00111010100000;     //80pi/512
   m_sin[81]  =  14'b11100101110001;     //81pi/512
   m_cos[81]  =  14'b00111010010111;     //81pi/512
   m_sin[82]  =  14'b11100101011101;     //82pi/512
   m_cos[82]  =  14'b00111010001111;     //82pi/512
   m_sin[83]  =  14'b11100101001010;     //83pi/512
   m_cos[83]  =  14'b00111010000110;     //83pi/512
   m_sin[84]  =  14'b11100100110110;     //84pi/512
   m_cos[84]  =  14'b00111001111101;     //84pi/512
   m_sin[85]  =  14'b11100100100011;     //85pi/512
   m_cos[85]  =  14'b00111001110100;     //85pi/512
   m_sin[86]  =  14'b11100100010000;     //86pi/512
   m_cos[86]  =  14'b00111001101010;     //86pi/512
   m_sin[87]  =  14'b11100011111101;     //87pi/512
   m_cos[87]  =  14'b00111001100001;     //87pi/512
   m_sin[88]  =  14'b11100011101001;     //88pi/512
   m_cos[88]  =  14'b00111001011000;     //88pi/512
   m_sin[89]  =  14'b11100011010110;     //89pi/512
   m_cos[89]  =  14'b00111001001110;     //89pi/512
   m_sin[90]  =  14'b11100011000011;     //90pi/512
   m_cos[90]  =  14'b00111001000100;     //90pi/512
   m_sin[91]  =  14'b11100010110000;     //91pi/512
   m_cos[91]  =  14'b00111000111011;     //91pi/512
   m_sin[92]  =  14'b11100010011101;     //92pi/512
   m_cos[92]  =  14'b00111000110001;     //92pi/512
   m_sin[93]  =  14'b11100010001010;     //93pi/512
   m_cos[93]  =  14'b00111000100111;     //93pi/512
   m_sin[94]  =  14'b11100001110111;     //94pi/512
   m_cos[94]  =  14'b00111000011101;     //94pi/512
   m_sin[95]  =  14'b11100001100101;     //95pi/512
   m_cos[95]  =  14'b00111000010011;     //95pi/512
   m_sin[96]  =  14'b11100001010010;     //96pi/512
   m_cos[96]  =  14'b00111000001001;     //96pi/512
   m_sin[97]  =  14'b11100000111111;     //97pi/512
   m_cos[97]  =  14'b00110111111110;     //97pi/512
   m_sin[98]  =  14'b11100000101100;     //98pi/512
   m_cos[98]  =  14'b00110111110100;     //98pi/512
   m_sin[99]  =  14'b11100000011010;     //99pi/512
   m_cos[99]  =  14'b00110111101010;     //99pi/512
   m_sin[100]  =  14'b11100000000111;     //100pi/512
   m_cos[100]  =  14'b00110111011111;     //100pi/512
   m_sin[101]  =  14'b11011111110101;     //101pi/512
   m_cos[101]  =  14'b00110111010100;     //101pi/512
   m_sin[102]  =  14'b11011111100010;     //102pi/512
   m_cos[102]  =  14'b00110111001001;     //102pi/512
   m_sin[103]  =  14'b11011111010000;     //103pi/512
   m_cos[103]  =  14'b00110110111111;     //103pi/512
   m_sin[104]  =  14'b11011110111110;     //104pi/512
   m_cos[104]  =  14'b00110110110100;     //104pi/512
   m_sin[105]  =  14'b11011110101011;     //105pi/512
   m_cos[105]  =  14'b00110110101001;     //105pi/512
   m_sin[106]  =  14'b11011110011001;     //106pi/512
   m_cos[106]  =  14'b00110110011101;     //106pi/512
   m_sin[107]  =  14'b11011110000111;     //107pi/512
   m_cos[107]  =  14'b00110110010010;     //107pi/512
   m_sin[108]  =  14'b11011101110101;     //108pi/512
   m_cos[108]  =  14'b00110110000111;     //108pi/512
   m_sin[109]  =  14'b11011101100011;     //109pi/512
   m_cos[109]  =  14'b00110101111011;     //109pi/512
   m_sin[110]  =  14'b11011101010001;     //110pi/512
   m_cos[110]  =  14'b00110101110000;     //110pi/512
   m_sin[111]  =  14'b11011100111111;     //111pi/512
   m_cos[111]  =  14'b00110101100100;     //111pi/512
   m_sin[112]  =  14'b11011100101101;     //112pi/512
   m_cos[112]  =  14'b00110101011000;     //112pi/512
   m_sin[113]  =  14'b11011100011011;     //113pi/512
   m_cos[113]  =  14'b00110101001101;     //113pi/512
   m_sin[114]  =  14'b11011100001010;     //114pi/512
   m_cos[114]  =  14'b00110101000001;     //114pi/512
   m_sin[115]  =  14'b11011011111000;     //115pi/512
   m_cos[115]  =  14'b00110100110101;     //115pi/512
   m_sin[116]  =  14'b11011011100110;     //116pi/512
   m_cos[116]  =  14'b00110100101000;     //116pi/512
   m_sin[117]  =  14'b11011011010101;     //117pi/512
   m_cos[117]  =  14'b00110100011100;     //117pi/512
   m_sin[118]  =  14'b11011011000011;     //118pi/512
   m_cos[118]  =  14'b00110100010000;     //118pi/512
   m_sin[119]  =  14'b11011010110010;     //119pi/512
   m_cos[119]  =  14'b00110100000100;     //119pi/512
   m_sin[120]  =  14'b11011010100001;     //120pi/512
   m_cos[120]  =  14'b00110011110111;     //120pi/512
   m_sin[121]  =  14'b11011010001111;     //121pi/512
   m_cos[121]  =  14'b00110011101011;     //121pi/512
   m_sin[122]  =  14'b11011001111110;     //122pi/512
   m_cos[122]  =  14'b00110011011110;     //122pi/512
   m_sin[123]  =  14'b11011001101101;     //123pi/512
   m_cos[123]  =  14'b00110011010001;     //123pi/512
   m_sin[124]  =  14'b11011001011100;     //124pi/512
   m_cos[124]  =  14'b00110011000100;     //124pi/512
   m_sin[125]  =  14'b11011001001011;     //125pi/512
   m_cos[125]  =  14'b00110010110111;     //125pi/512
   m_sin[126]  =  14'b11011000111010;     //126pi/512
   m_cos[126]  =  14'b00110010101010;     //126pi/512
   m_sin[127]  =  14'b11011000101001;     //127pi/512
   m_cos[127]  =  14'b00110010011101;     //127pi/512
   m_sin[128]  =  14'b11011000011000;     //128pi/512
   m_cos[128]  =  14'b00110010010000;     //128pi/512
   m_sin[129]  =  14'b11011000000111;     //129pi/512
   m_cos[129]  =  14'b00110010000011;     //129pi/512
   m_sin[130]  =  14'b11010111110111;     //130pi/512
   m_cos[130]  =  14'b00110001110110;     //130pi/512
   m_sin[131]  =  14'b11010111100110;     //131pi/512
   m_cos[131]  =  14'b00110001101000;     //131pi/512
   m_sin[132]  =  14'b11010111010110;     //132pi/512
   m_cos[132]  =  14'b00110001011011;     //132pi/512
   m_sin[133]  =  14'b11010111000101;     //133pi/512
   m_cos[133]  =  14'b00110001001101;     //133pi/512
   m_sin[134]  =  14'b11010110110101;     //134pi/512
   m_cos[134]  =  14'b00110000111111;     //134pi/512
   m_sin[135]  =  14'b11010110100100;     //135pi/512
   m_cos[135]  =  14'b00110000110001;     //135pi/512
   m_sin[136]  =  14'b11010110010100;     //136pi/512
   m_cos[136]  =  14'b00110000100100;     //136pi/512
   m_sin[137]  =  14'b11010110000100;     //137pi/512
   m_cos[137]  =  14'b00110000010110;     //137pi/512
   m_sin[138]  =  14'b11010101110100;     //138pi/512
   m_cos[138]  =  14'b00110000001000;     //138pi/512
   m_sin[139]  =  14'b11010101100100;     //139pi/512
   m_cos[139]  =  14'b00101111111001;     //139pi/512
   m_sin[140]  =  14'b11010101010100;     //140pi/512
   m_cos[140]  =  14'b00101111101011;     //140pi/512
   m_sin[141]  =  14'b11010101000100;     //141pi/512
   m_cos[141]  =  14'b00101111011101;     //141pi/512
   m_sin[142]  =  14'b11010100110100;     //142pi/512
   m_cos[142]  =  14'b00101111001111;     //142pi/512
   m_sin[143]  =  14'b11010100100101;     //143pi/512
   m_cos[143]  =  14'b00101111000000;     //143pi/512
   m_sin[144]  =  14'b11010100010101;     //144pi/512
   m_cos[144]  =  14'b00101110110010;     //144pi/512
   m_sin[145]  =  14'b11010100000101;     //145pi/512
   m_cos[145]  =  14'b00101110100011;     //145pi/512
   m_sin[146]  =  14'b11010011110110;     //146pi/512
   m_cos[146]  =  14'b00101110010100;     //146pi/512
   m_sin[147]  =  14'b11010011100110;     //147pi/512
   m_cos[147]  =  14'b00101110000110;     //147pi/512
   m_sin[148]  =  14'b11010011010111;     //148pi/512
   m_cos[148]  =  14'b00101101110111;     //148pi/512
   m_sin[149]  =  14'b11010011001000;     //149pi/512
   m_cos[149]  =  14'b00101101101000;     //149pi/512
   m_sin[150]  =  14'b11010010111001;     //150pi/512
   m_cos[150]  =  14'b00101101011001;     //150pi/512
   m_sin[151]  =  14'b11010010101001;     //151pi/512
   m_cos[151]  =  14'b00101101001010;     //151pi/512
   m_sin[152]  =  14'b11010010011010;     //152pi/512
   m_cos[152]  =  14'b00101100111010;     //152pi/512
   m_sin[153]  =  14'b11010010001011;     //153pi/512
   m_cos[153]  =  14'b00101100101011;     //153pi/512
   m_sin[154]  =  14'b11010001111101;     //154pi/512
   m_cos[154]  =  14'b00101100011100;     //154pi/512
   m_sin[155]  =  14'b11010001101110;     //155pi/512
   m_cos[155]  =  14'b00101100001100;     //155pi/512
   m_sin[156]  =  14'b11010001011111;     //156pi/512
   m_cos[156]  =  14'b00101011111101;     //156pi/512
   m_sin[157]  =  14'b11010001010000;     //157pi/512
   m_cos[157]  =  14'b00101011101101;     //157pi/512
   m_sin[158]  =  14'b11010001000010;     //158pi/512
   m_cos[158]  =  14'b00101011011110;     //158pi/512
   m_sin[159]  =  14'b11010000110011;     //159pi/512
   m_cos[159]  =  14'b00101011001110;     //159pi/512
   m_sin[160]  =  14'b11010000100101;     //160pi/512
   m_cos[160]  =  14'b00101010111110;     //160pi/512
   m_sin[161]  =  14'b11010000010111;     //161pi/512
   m_cos[161]  =  14'b00101010101110;     //161pi/512
   m_sin[162]  =  14'b11010000001001;     //162pi/512
   m_cos[162]  =  14'b00101010011110;     //162pi/512
   m_sin[163]  =  14'b11001111111010;     //163pi/512
   m_cos[163]  =  14'b00101010001110;     //163pi/512
   m_sin[164]  =  14'b11001111101100;     //164pi/512
   m_cos[164]  =  14'b00101001111110;     //164pi/512
   m_sin[165]  =  14'b11001111011110;     //165pi/512
   m_cos[165]  =  14'b00101001101110;     //165pi/512
   m_sin[166]  =  14'b11001111010000;     //166pi/512
   m_cos[166]  =  14'b00101001011110;     //166pi/512
   m_sin[167]  =  14'b11001111000011;     //167pi/512
   m_cos[167]  =  14'b00101001001110;     //167pi/512
   m_sin[168]  =  14'b11001110110101;     //168pi/512
   m_cos[168]  =  14'b00101000111101;     //168pi/512
   m_sin[169]  =  14'b11001110100111;     //169pi/512
   m_cos[169]  =  14'b00101000101101;     //169pi/512
   m_sin[170]  =  14'b11001110011010;     //170pi/512
   m_cos[170]  =  14'b00101000011100;     //170pi/512
   m_sin[171]  =  14'b11001110001100;     //171pi/512
   m_cos[171]  =  14'b00101000001100;     //171pi/512
   m_sin[172]  =  14'b11001101111111;     //172pi/512
   m_cos[172]  =  14'b00100111111011;     //172pi/512
   m_sin[173]  =  14'b11001101110010;     //173pi/512
   m_cos[173]  =  14'b00100111101010;     //173pi/512
   m_sin[174]  =  14'b11001101100100;     //174pi/512
   m_cos[174]  =  14'b00100111011001;     //174pi/512
   m_sin[175]  =  14'b11001101010111;     //175pi/512
   m_cos[175]  =  14'b00100111001001;     //175pi/512
   m_sin[176]  =  14'b11001101001010;     //176pi/512
   m_cos[176]  =  14'b00100110111000;     //176pi/512
   m_sin[177]  =  14'b11001100111101;     //177pi/512
   m_cos[177]  =  14'b00100110100111;     //177pi/512
   m_sin[178]  =  14'b11001100110001;     //178pi/512
   m_cos[178]  =  14'b00100110010110;     //178pi/512
   m_sin[179]  =  14'b11001100100100;     //179pi/512
   m_cos[179]  =  14'b00100110000100;     //179pi/512
   m_sin[180]  =  14'b11001100010111;     //180pi/512
   m_cos[180]  =  14'b00100101110011;     //180pi/512
   m_sin[181]  =  14'b11001100001011;     //181pi/512
   m_cos[181]  =  14'b00100101100010;     //181pi/512
   m_sin[182]  =  14'b11001011111110;     //182pi/512
   m_cos[182]  =  14'b00100101010001;     //182pi/512
   m_sin[183]  =  14'b11001011110010;     //183pi/512
   m_cos[183]  =  14'b00100100111111;     //183pi/512
   m_sin[184]  =  14'b11001011100101;     //184pi/512
   m_cos[184]  =  14'b00100100101110;     //184pi/512
   m_sin[185]  =  14'b11001011011001;     //185pi/512
   m_cos[185]  =  14'b00100100011100;     //185pi/512
   m_sin[186]  =  14'b11001011001101;     //186pi/512
   m_cos[186]  =  14'b00100100001011;     //186pi/512
   m_sin[187]  =  14'b11001011000001;     //187pi/512
   m_cos[187]  =  14'b00100011111001;     //187pi/512
   m_sin[188]  =  14'b11001010110101;     //188pi/512
   m_cos[188]  =  14'b00100011100111;     //188pi/512
   m_sin[189]  =  14'b11001010101001;     //189pi/512
   m_cos[189]  =  14'b00100011010110;     //189pi/512
   m_sin[190]  =  14'b11001010011110;     //190pi/512
   m_cos[190]  =  14'b00100011000100;     //190pi/512
   m_sin[191]  =  14'b11001010010010;     //191pi/512
   m_cos[191]  =  14'b00100010110010;     //191pi/512
   m_sin[192]  =  14'b11001010000110;     //192pi/512
   m_cos[192]  =  14'b00100010100000;     //192pi/512
   m_sin[193]  =  14'b11001001111011;     //193pi/512
   m_cos[193]  =  14'b00100010001110;     //193pi/512
   m_sin[194]  =  14'b11001001101111;     //194pi/512
   m_cos[194]  =  14'b00100001111100;     //194pi/512
   m_sin[195]  =  14'b11001001100100;     //195pi/512
   m_cos[195]  =  14'b00100001101010;     //195pi/512
   m_sin[196]  =  14'b11001001011001;     //196pi/512
   m_cos[196]  =  14'b00100001010111;     //196pi/512
   m_sin[197]  =  14'b11001001001110;     //197pi/512
   m_cos[197]  =  14'b00100001000101;     //197pi/512
   m_sin[198]  =  14'b11001001000011;     //198pi/512
   m_cos[198]  =  14'b00100000110011;     //198pi/512
   m_sin[199]  =  14'b11001000111000;     //199pi/512
   m_cos[199]  =  14'b00100000100000;     //199pi/512
   m_sin[200]  =  14'b11001000101101;     //200pi/512
   m_cos[200]  =  14'b00100000001110;     //200pi/512
   m_sin[201]  =  14'b11001000100010;     //201pi/512
   m_cos[201]  =  14'b00011111111100;     //201pi/512
   m_sin[202]  =  14'b11001000011000;     //202pi/512
   m_cos[202]  =  14'b00011111101001;     //202pi/512
   m_sin[203]  =  14'b11001000001101;     //203pi/512
   m_cos[203]  =  14'b00011111010110;     //203pi/512
   m_sin[204]  =  14'b11001000000011;     //204pi/512
   m_cos[204]  =  14'b00011111000100;     //204pi/512
   m_sin[205]  =  14'b11000111111001;     //205pi/512
   m_cos[205]  =  14'b00011110110001;     //205pi/512
   m_sin[206]  =  14'b11000111101110;     //206pi/512
   m_cos[206]  =  14'b00011110011110;     //206pi/512
   m_sin[207]  =  14'b11000111100100;     //207pi/512
   m_cos[207]  =  14'b00011110001011;     //207pi/512
   m_sin[208]  =  14'b11000111011010;     //208pi/512
   m_cos[208]  =  14'b00011101111001;     //208pi/512
   m_sin[209]  =  14'b11000111010000;     //209pi/512
   m_cos[209]  =  14'b00011101100110;     //209pi/512
   m_sin[210]  =  14'b11000111000110;     //210pi/512
   m_cos[210]  =  14'b00011101010011;     //210pi/512
   m_sin[211]  =  14'b11000110111101;     //211pi/512
   m_cos[211]  =  14'b00011101000000;     //211pi/512
   m_sin[212]  =  14'b11000110110011;     //212pi/512
   m_cos[212]  =  14'b00011100101101;     //212pi/512
   m_sin[213]  =  14'b11000110101010;     //213pi/512
   m_cos[213]  =  14'b00011100011001;     //213pi/512
   m_sin[214]  =  14'b11000110100000;     //214pi/512
   m_cos[214]  =  14'b00011100000110;     //214pi/512
   m_sin[215]  =  14'b11000110010111;     //215pi/512
   m_cos[215]  =  14'b00011011110011;     //215pi/512
   m_sin[216]  =  14'b11000110001110;     //216pi/512
   m_cos[216]  =  14'b00011011100000;     //216pi/512
   m_sin[217]  =  14'b11000110000100;     //217pi/512
   m_cos[217]  =  14'b00011011001101;     //217pi/512
   m_sin[218]  =  14'b11000101111011;     //218pi/512
   m_cos[218]  =  14'b00011010111001;     //218pi/512
   m_sin[219]  =  14'b11000101110010;     //219pi/512
   m_cos[219]  =  14'b00011010100110;     //219pi/512
   m_sin[220]  =  14'b11000101101010;     //220pi/512
   m_cos[220]  =  14'b00011010010010;     //220pi/512
   m_sin[221]  =  14'b11000101100001;     //221pi/512
   m_cos[221]  =  14'b00011001111111;     //221pi/512
   m_sin[222]  =  14'b11000101011000;     //222pi/512
   m_cos[222]  =  14'b00011001101011;     //222pi/512
   m_sin[223]  =  14'b11000101010000;     //223pi/512
   m_cos[223]  =  14'b00011001011000;     //223pi/512
   m_sin[224]  =  14'b11000101000111;     //224pi/512
   m_cos[224]  =  14'b00011001000100;     //224pi/512
   m_sin[225]  =  14'b11000100111111;     //225pi/512
   m_cos[225]  =  14'b00011000110000;     //225pi/512
   m_sin[226]  =  14'b11000100110111;     //226pi/512
   m_cos[226]  =  14'b00011000011101;     //226pi/512
   m_sin[227]  =  14'b11000100101111;     //227pi/512
   m_cos[227]  =  14'b00011000001001;     //227pi/512
   m_sin[228]  =  14'b11000100100111;     //228pi/512
   m_cos[228]  =  14'b00010111110101;     //228pi/512
   m_sin[229]  =  14'b11000100011111;     //229pi/512
   m_cos[229]  =  14'b00010111100001;     //229pi/512
   m_sin[230]  =  14'b11000100010111;     //230pi/512
   m_cos[230]  =  14'b00010111001101;     //230pi/512
   m_sin[231]  =  14'b11000100001111;     //231pi/512
   m_cos[231]  =  14'b00010110111001;     //231pi/512
   m_sin[232]  =  14'b11000100001000;     //232pi/512
   m_cos[232]  =  14'b00010110100101;     //232pi/512
   m_sin[233]  =  14'b11000100000000;     //233pi/512
   m_cos[233]  =  14'b00010110010001;     //233pi/512
   m_sin[234]  =  14'b11000011111001;     //234pi/512
   m_cos[234]  =  14'b00010101111101;     //234pi/512
   m_sin[235]  =  14'b11000011110010;     //235pi/512
   m_cos[235]  =  14'b00010101101001;     //235pi/512
   m_sin[236]  =  14'b11000011101010;     //236pi/512
   m_cos[236]  =  14'b00010101010101;     //236pi/512
   m_sin[237]  =  14'b11000011100011;     //237pi/512
   m_cos[237]  =  14'b00010101000001;     //237pi/512
   m_sin[238]  =  14'b11000011011100;     //238pi/512
   m_cos[238]  =  14'b00010100101101;     //238pi/512
   m_sin[239]  =  14'b11000011010101;     //239pi/512
   m_cos[239]  =  14'b00010100011001;     //239pi/512
   m_sin[240]  =  14'b11000011001111;     //240pi/512
   m_cos[240]  =  14'b00010100000100;     //240pi/512
   m_sin[241]  =  14'b11000011001000;     //241pi/512
   m_cos[241]  =  14'b00010011110000;     //241pi/512
   m_sin[242]  =  14'b11000011000010;     //242pi/512
   m_cos[242]  =  14'b00010011011100;     //242pi/512
   m_sin[243]  =  14'b11000010111011;     //243pi/512
   m_cos[243]  =  14'b00010011000111;     //243pi/512
   m_sin[244]  =  14'b11000010110101;     //244pi/512
   m_cos[244]  =  14'b00010010110011;     //244pi/512
   m_sin[245]  =  14'b11000010101111;     //245pi/512
   m_cos[245]  =  14'b00010010011110;     //245pi/512
   m_sin[246]  =  14'b11000010101000;     //246pi/512
   m_cos[246]  =  14'b00010010001010;     //246pi/512
   m_sin[247]  =  14'b11000010100010;     //247pi/512
   m_cos[247]  =  14'b00010001110110;     //247pi/512
   m_sin[248]  =  14'b11000010011101;     //248pi/512
   m_cos[248]  =  14'b00010001100001;     //248pi/512
   m_sin[249]  =  14'b11000010010111;     //249pi/512
   m_cos[249]  =  14'b00010001001100;     //249pi/512
   m_sin[250]  =  14'b11000010010001;     //250pi/512
   m_cos[250]  =  14'b00010000111000;     //250pi/512
   m_sin[251]  =  14'b11000010001011;     //251pi/512
   m_cos[251]  =  14'b00010000100011;     //251pi/512
   m_sin[252]  =  14'b11000010000110;     //252pi/512
   m_cos[252]  =  14'b00010000001111;     //252pi/512
   m_sin[253]  =  14'b11000010000001;     //253pi/512
   m_cos[253]  =  14'b00001111111010;     //253pi/512
   m_sin[254]  =  14'b11000001111011;     //254pi/512
   m_cos[254]  =  14'b00001111100101;     //254pi/512
   m_sin[255]  =  14'b11000001110110;     //255pi/512
   m_cos[255]  =  14'b00001111010000;     //255pi/512
   m_sin[256]  =  14'b11000001110001;     //256pi/512
   m_cos[256]  =  14'b00001110111100;     //256pi/512
   m_sin[257]  =  14'b11000001101100;     //257pi/512
   m_cos[257]  =  14'b00001110100111;     //257pi/512
   m_sin[258]  =  14'b11000001100111;     //258pi/512
   m_cos[258]  =  14'b00001110010010;     //258pi/512
   m_sin[259]  =  14'b11000001100011;     //259pi/512
   m_cos[259]  =  14'b00001101111101;     //259pi/512
   m_sin[260]  =  14'b11000001011110;     //260pi/512
   m_cos[260]  =  14'b00001101101000;     //260pi/512
   m_sin[261]  =  14'b11000001011010;     //261pi/512
   m_cos[261]  =  14'b00001101010100;     //261pi/512
   m_sin[262]  =  14'b11000001010101;     //262pi/512
   m_cos[262]  =  14'b00001100111111;     //262pi/512
   m_sin[263]  =  14'b11000001010001;     //263pi/512
   m_cos[263]  =  14'b00001100101010;     //263pi/512
   m_sin[264]  =  14'b11000001001101;     //264pi/512
   m_cos[264]  =  14'b00001100010101;     //264pi/512
   m_sin[265]  =  14'b11000001001001;     //265pi/512
   m_cos[265]  =  14'b00001100000000;     //265pi/512
   m_sin[266]  =  14'b11000001000101;     //266pi/512
   m_cos[266]  =  14'b00001011101011;     //266pi/512
   m_sin[267]  =  14'b11000001000001;     //267pi/512
   m_cos[267]  =  14'b00001011010110;     //267pi/512
   m_sin[268]  =  14'b11000000111101;     //268pi/512
   m_cos[268]  =  14'b00001011000001;     //268pi/512
   m_sin[269]  =  14'b11000000111010;     //269pi/512
   m_cos[269]  =  14'b00001010101100;     //269pi/512
   m_sin[270]  =  14'b11000000110110;     //270pi/512
   m_cos[270]  =  14'b00001010010111;     //270pi/512
   m_sin[271]  =  14'b11000000110011;     //271pi/512
   m_cos[271]  =  14'b00001010000001;     //271pi/512
   m_sin[272]  =  14'b11000000101111;     //272pi/512
   m_cos[272]  =  14'b00001001101100;     //272pi/512
   m_sin[273]  =  14'b11000000101100;     //273pi/512
   m_cos[273]  =  14'b00001001010111;     //273pi/512
   m_sin[274]  =  14'b11000000101001;     //274pi/512
   m_cos[274]  =  14'b00001001000010;     //274pi/512
   m_sin[275]  =  14'b11000000100110;     //275pi/512
   m_cos[275]  =  14'b00001000101101;     //275pi/512
   m_sin[276]  =  14'b11000000100011;     //276pi/512
   m_cos[276]  =  14'b00001000011000;     //276pi/512
   m_sin[277]  =  14'b11000000100001;     //277pi/512
   m_cos[277]  =  14'b00001000000011;     //277pi/512
   m_sin[278]  =  14'b11000000011110;     //278pi/512
   m_cos[278]  =  14'b00000111101101;     //278pi/512
   m_sin[279]  =  14'b11000000011011;     //279pi/512
   m_cos[279]  =  14'b00000111011000;     //279pi/512
   m_sin[280]  =  14'b11000000011001;     //280pi/512
   m_cos[280]  =  14'b00000111000011;     //280pi/512
   m_sin[281]  =  14'b11000000010111;     //281pi/512
   m_cos[281]  =  14'b00000110101110;     //281pi/512
   m_sin[282]  =  14'b11000000010100;     //282pi/512
   m_cos[282]  =  14'b00000110011000;     //282pi/512
   m_sin[283]  =  14'b11000000010010;     //283pi/512
   m_cos[283]  =  14'b00000110000011;     //283pi/512
   m_sin[284]  =  14'b11000000010000;     //284pi/512
   m_cos[284]  =  14'b00000101101110;     //284pi/512
   m_sin[285]  =  14'b11000000001111;     //285pi/512
   m_cos[285]  =  14'b00000101011001;     //285pi/512
   m_sin[286]  =  14'b11000000001101;     //286pi/512
   m_cos[286]  =  14'b00000101000011;     //286pi/512
   m_sin[287]  =  14'b11000000001011;     //287pi/512
   m_cos[287]  =  14'b00000100101110;     //287pi/512
   m_sin[288]  =  14'b11000000001010;     //288pi/512
   m_cos[288]  =  14'b00000100011001;     //288pi/512
   m_sin[289]  =  14'b11000000001000;     //289pi/512
   m_cos[289]  =  14'b00000100000011;     //289pi/512
   m_sin[290]  =  14'b11000000000111;     //290pi/512
   m_cos[290]  =  14'b00000011101110;     //290pi/512
   m_sin[291]  =  14'b11000000000110;     //291pi/512
   m_cos[291]  =  14'b00000011011001;     //291pi/512
   m_sin[292]  =  14'b11000000000101;     //292pi/512
   m_cos[292]  =  14'b00000011000011;     //292pi/512
   m_sin[293]  =  14'b11000000000100;     //293pi/512
   m_cos[293]  =  14'b00000010101110;     //293pi/512
   m_sin[294]  =  14'b11000000000011;     //294pi/512
   m_cos[294]  =  14'b00000010011001;     //294pi/512
   m_sin[295]  =  14'b11000000000010;     //295pi/512
   m_cos[295]  =  14'b00000010000011;     //295pi/512
   m_sin[296]  =  14'b11000000000001;     //296pi/512
   m_cos[296]  =  14'b00000001101110;     //296pi/512
   m_sin[297]  =  14'b11000000000001;     //297pi/512
   m_cos[297]  =  14'b00000001011001;     //297pi/512
   m_sin[298]  =  14'b11000000000001;     //298pi/512
   m_cos[298]  =  14'b00000001000011;     //298pi/512
   m_sin[299]  =  14'b11000000000000;     //299pi/512
   m_cos[299]  =  14'b00000000101110;     //299pi/512
   m_sin[300]  =  14'b11000000000000;     //300pi/512
   m_cos[300]  =  14'b00000000011001;     //300pi/512
   m_sin[301]  =  14'b11000000000000;     //301pi/512
   m_cos[301]  =  14'b00000000000011;     //301pi/512
   m_sin[302]  =  14'b11000000000000;     //302pi/512
   m_cos[302]  =  14'b11111111101110;     //302pi/512
   m_sin[303]  =  14'b11000000000000;     //303pi/512
   m_cos[303]  =  14'b11111111011001;     //303pi/512
   m_sin[304]  =  14'b11000000000000;     //304pi/512
   m_cos[304]  =  14'b11111111000100;     //304pi/512
   m_sin[305]  =  14'b11000000000001;     //305pi/512
   m_cos[305]  =  14'b11111110101110;     //305pi/512
   m_sin[306]  =  14'b11000000000001;     //306pi/512
   m_cos[306]  =  14'b11111110011001;     //306pi/512
   m_sin[307]  =  14'b11000000000010;     //307pi/512
   m_cos[307]  =  14'b11111110000100;     //307pi/512
   m_sin[308]  =  14'b11000000000011;     //308pi/512
   m_cos[308]  =  14'b11111101101110;     //308pi/512
   m_sin[309]  =  14'b11000000000011;     //309pi/512
   m_cos[309]  =  14'b11111101011001;     //309pi/512
   m_sin[310]  =  14'b11000000000100;     //310pi/512
   m_cos[310]  =  14'b11111101000100;     //310pi/512
   m_sin[311]  =  14'b11000000000101;     //311pi/512
   m_cos[311]  =  14'b11111100101110;     //311pi/512
   m_sin[312]  =  14'b11000000000111;     //312pi/512
   m_cos[312]  =  14'b11111100011001;     //312pi/512
   m_sin[313]  =  14'b11000000001000;     //313pi/512
   m_cos[313]  =  14'b11111100000100;     //313pi/512
   m_sin[314]  =  14'b11000000001001;     //314pi/512
   m_cos[314]  =  14'b11111011101110;     //314pi/512
   m_sin[315]  =  14'b11000000001011;     //315pi/512
   m_cos[315]  =  14'b11111011011001;     //315pi/512
   m_sin[316]  =  14'b11000000001100;     //316pi/512
   m_cos[316]  =  14'b11111011000100;     //316pi/512
   m_sin[317]  =  14'b11000000001110;     //317pi/512
   m_cos[317]  =  14'b11111010101110;     //317pi/512
   m_sin[318]  =  14'b11000000010000;     //318pi/512
   m_cos[318]  =  14'b11111010011001;     //318pi/512
   m_sin[319]  =  14'b11000000010010;     //319pi/512
   m_cos[319]  =  14'b11111010000100;     //319pi/512
   m_sin[320]  =  14'b11000000010100;     //320pi/512
   m_cos[320]  =  14'b11111001101111;     //320pi/512
   m_sin[321]  =  14'b11000000010110;     //321pi/512
   m_cos[321]  =  14'b11111001011001;     //321pi/512
   m_sin[322]  =  14'b11000000011000;     //322pi/512
   m_cos[322]  =  14'b11111001000100;     //322pi/512
   m_sin[323]  =  14'b11000000011011;     //323pi/512
   m_cos[323]  =  14'b11111000101111;     //323pi/512
   m_sin[324]  =  14'b11000000011101;     //324pi/512
   m_cos[324]  =  14'b11111000011010;     //324pi/512
   m_sin[325]  =  14'b11000000100000;     //325pi/512
   m_cos[325]  =  14'b11111000000100;     //325pi/512
   m_sin[326]  =  14'b11000000100010;     //326pi/512
   m_cos[326]  =  14'b11110111101111;     //326pi/512
   m_sin[327]  =  14'b11000000100101;     //327pi/512
   m_cos[327]  =  14'b11110111011010;     //327pi/512
   m_sin[328]  =  14'b11000000101000;     //328pi/512
   m_cos[328]  =  14'b11110111000101;     //328pi/512
   m_sin[329]  =  14'b11000000101011;     //329pi/512
   m_cos[329]  =  14'b11110110110000;     //329pi/512
   m_sin[330]  =  14'b11000000101110;     //330pi/512
   m_cos[330]  =  14'b11110110011011;     //330pi/512
   m_sin[331]  =  14'b11000000110001;     //331pi/512
   m_cos[331]  =  14'b11110110000101;     //331pi/512
   m_sin[332]  =  14'b11000000110101;     //332pi/512
   m_cos[332]  =  14'b11110101110000;     //332pi/512
   m_sin[333]  =  14'b11000000111000;     //333pi/512
   m_cos[333]  =  14'b11110101011011;     //333pi/512
   m_sin[334]  =  14'b11000000111100;     //334pi/512
   m_cos[334]  =  14'b11110101000110;     //334pi/512
   m_sin[335]  =  14'b11000001000000;     //335pi/512
   m_cos[335]  =  14'b11110100110001;     //335pi/512
   m_sin[336]  =  14'b11000001000011;     //336pi/512
   m_cos[336]  =  14'b11110100011100;     //336pi/512
   m_sin[337]  =  14'b11000001000111;     //337pi/512
   m_cos[337]  =  14'b11110100000111;     //337pi/512
   m_sin[338]  =  14'b11000001001011;     //338pi/512
   m_cos[338]  =  14'b11110011110010;     //338pi/512
   m_sin[339]  =  14'b11000001001111;     //339pi/512
   m_cos[339]  =  14'b11110011011101;     //339pi/512
   m_sin[340]  =  14'b11000001010100;     //340pi/512
   m_cos[340]  =  14'b11110011001000;     //340pi/512
   m_sin[341]  =  14'b11000001011000;     //341pi/512
   m_cos[341]  =  14'b11110010110011;     //341pi/512
   m_sin[342]  =  14'b11000001011100;     //342pi/512
   m_cos[342]  =  14'b11110010011110;     //342pi/512
   m_sin[343]  =  14'b11000001100001;     //343pi/512
   m_cos[343]  =  14'b11110010001010;     //343pi/512
   m_sin[344]  =  14'b11000001100110;     //344pi/512
   m_cos[344]  =  14'b11110001110101;     //344pi/512
   m_sin[345]  =  14'b11000001101011;     //345pi/512
   m_cos[345]  =  14'b11110001100000;     //345pi/512
   m_sin[346]  =  14'b11000001101111;     //346pi/512
   m_cos[346]  =  14'b11110001001011;     //346pi/512
   m_sin[347]  =  14'b11000001110100;     //347pi/512
   m_cos[347]  =  14'b11110000110110;     //347pi/512
   m_sin[348]  =  14'b11000001111010;     //348pi/512
   m_cos[348]  =  14'b11110000100010;     //348pi/512
   m_sin[349]  =  14'b11000001111111;     //349pi/512
   m_cos[349]  =  14'b11110000001101;     //349pi/512
   m_sin[350]  =  14'b11000010000100;     //350pi/512
   m_cos[350]  =  14'b11101111111000;     //350pi/512
   m_sin[351]  =  14'b11000010001010;     //351pi/512
   m_cos[351]  =  14'b11101111100100;     //351pi/512
   m_sin[352]  =  14'b11000010001111;     //352pi/512
   m_cos[352]  =  14'b11101111001111;     //352pi/512
   m_sin[353]  =  14'b11000010010101;     //353pi/512
   m_cos[353]  =  14'b11101110111010;     //353pi/512
   m_sin[354]  =  14'b11000010011010;     //354pi/512
   m_cos[354]  =  14'b11101110100110;     //354pi/512
   m_sin[355]  =  14'b11000010100000;     //355pi/512
   m_cos[355]  =  14'b11101110010001;     //355pi/512
   m_sin[356]  =  14'b11000010100110;     //356pi/512
   m_cos[356]  =  14'b11101101111101;     //356pi/512
   m_sin[357]  =  14'b11000010101100;     //357pi/512
   m_cos[357]  =  14'b11101101101000;     //357pi/512
   m_sin[358]  =  14'b11000010110011;     //358pi/512
   m_cos[358]  =  14'b11101101010100;     //358pi/512
   m_sin[359]  =  14'b11000010111001;     //359pi/512
   m_cos[359]  =  14'b11101100111111;     //359pi/512
   m_sin[360]  =  14'b11000010111111;     //360pi/512
   m_cos[360]  =  14'b11101100101011;     //360pi/512
   m_sin[361]  =  14'b11000011000110;     //361pi/512
   m_cos[361]  =  14'b11101100010111;     //361pi/512
   m_sin[362]  =  14'b11000011001100;     //362pi/512
   m_cos[362]  =  14'b11101100000010;     //362pi/512
   m_sin[363]  =  14'b11000011010011;     //363pi/512
   m_cos[363]  =  14'b11101011101110;     //363pi/512
   m_sin[364]  =  14'b11000011011010;     //364pi/512
   m_cos[364]  =  14'b11101011011010;     //364pi/512
   m_sin[365]  =  14'b11000011100001;     //365pi/512
   m_cos[365]  =  14'b11101011000110;     //365pi/512
   m_sin[366]  =  14'b11000011101000;     //366pi/512
   m_cos[366]  =  14'b11101010110001;     //366pi/512
   m_sin[367]  =  14'b11000011101111;     //367pi/512
   m_cos[367]  =  14'b11101010011101;     //367pi/512
   m_sin[368]  =  14'b11000011110110;     //368pi/512
   m_cos[368]  =  14'b11101010001001;     //368pi/512
   m_sin[369]  =  14'b11000011111110;     //369pi/512
   m_cos[369]  =  14'b11101001110101;     //369pi/512
   m_sin[370]  =  14'b11000100000101;     //370pi/512
   m_cos[370]  =  14'b11101001100001;     //370pi/512
   m_sin[371]  =  14'b11000100001101;     //371pi/512
   m_cos[371]  =  14'b11101001001101;     //371pi/512
   m_sin[372]  =  14'b11000100010100;     //372pi/512
   m_cos[372]  =  14'b11101000111001;     //372pi/512
   m_sin[373]  =  14'b11000100011100;     //373pi/512
   m_cos[373]  =  14'b11101000100101;     //373pi/512
   m_sin[374]  =  14'b11000100100100;     //374pi/512
   m_cos[374]  =  14'b11101000010001;     //374pi/512
   m_sin[375]  =  14'b11000100101100;     //375pi/512
   m_cos[375]  =  14'b11100111111110;     //375pi/512
   m_sin[376]  =  14'b11000100110100;     //376pi/512
   m_cos[376]  =  14'b11100111101010;     //376pi/512
   m_sin[377]  =  14'b11000100111100;     //377pi/512
   m_cos[377]  =  14'b11100111010110;     //377pi/512
   m_sin[378]  =  14'b11000101000100;     //378pi/512
   m_cos[378]  =  14'b11100111000010;     //378pi/512
   m_sin[379]  =  14'b11000101001101;     //379pi/512
   m_cos[379]  =  14'b11100110101111;     //379pi/512
   m_sin[380]  =  14'b11000101010101;     //380pi/512
   m_cos[380]  =  14'b11100110011011;     //380pi/512
   m_sin[381]  =  14'b11000101011110;     //381pi/512
   m_cos[381]  =  14'b11100110001000;     //381pi/512
   m_sin[382]  =  14'b11000101100111;     //382pi/512
   m_cos[382]  =  14'b11100101110100;     //382pi/512
   m_sin[383]  =  14'b11000101101111;     //383pi/512
   m_cos[383]  =  14'b11100101100001;     //383pi/512
   m_sin[384]  =  14'b11000101111000;     //384pi/512
   m_cos[384]  =  14'b11100101001101;     //384pi/512
   m_sin[385]  =  14'b11000110000001;     //385pi/512
   m_cos[385]  =  14'b11100100111010;     //385pi/512
   m_sin[386]  =  14'b11000110001010;     //386pi/512
   m_cos[386]  =  14'b11100100100110;     //386pi/512
   m_sin[387]  =  14'b11000110010100;     //387pi/512
   m_cos[387]  =  14'b11100100010011;     //387pi/512
   m_sin[388]  =  14'b11000110011101;     //388pi/512
   m_cos[388]  =  14'b11100100000000;     //388pi/512
   m_sin[389]  =  14'b11000110100110;     //389pi/512
   m_cos[389]  =  14'b11100011101101;     //389pi/512
   m_sin[390]  =  14'b11000110110000;     //390pi/512
   m_cos[390]  =  14'b11100011011010;     //390pi/512
   m_sin[391]  =  14'b11000110111001;     //391pi/512
   m_cos[391]  =  14'b11100011000111;     //391pi/512
   m_sin[392]  =  14'b11000111000011;     //392pi/512
   m_cos[392]  =  14'b11100010110100;     //392pi/512
   m_sin[393]  =  14'b11000111001101;     //393pi/512
   m_cos[393]  =  14'b11100010100001;     //393pi/512
   m_sin[394]  =  14'b11000111010111;     //394pi/512
   m_cos[394]  =  14'b11100010001110;     //394pi/512
   m_sin[395]  =  14'b11000111100001;     //395pi/512
   m_cos[395]  =  14'b11100001111011;     //395pi/512
   m_sin[396]  =  14'b11000111101011;     //396pi/512
   m_cos[396]  =  14'b11100001101000;     //396pi/512
   m_sin[397]  =  14'b11000111110101;     //397pi/512
   m_cos[397]  =  14'b11100001010101;     //397pi/512
   m_sin[398]  =  14'b11000111111111;     //398pi/512
   m_cos[398]  =  14'b11100001000010;     //398pi/512
   m_sin[399]  =  14'b11001000001010;     //399pi/512
   m_cos[399]  =  14'b11100000110000;     //399pi/512
   m_sin[400]  =  14'b11001000010100;     //400pi/512
   m_cos[400]  =  14'b11100000011101;     //400pi/512
   m_sin[401]  =  14'b11001000011111;     //401pi/512
   m_cos[401]  =  14'b11100000001011;     //401pi/512
   m_sin[402]  =  14'b11001000101001;     //402pi/512
   m_cos[402]  =  14'b11011111111000;     //402pi/512
   m_sin[403]  =  14'b11001000110100;     //403pi/512
   m_cos[403]  =  14'b11011111100110;     //403pi/512
   m_sin[404]  =  14'b11001000111111;     //404pi/512
   m_cos[404]  =  14'b11011111010011;     //404pi/512
   m_sin[405]  =  14'b11001001001010;     //405pi/512
   m_cos[405]  =  14'b11011111000001;     //405pi/512
   m_sin[406]  =  14'b11001001010101;     //406pi/512
   m_cos[406]  =  14'b11011110101111;     //406pi/512
   m_sin[407]  =  14'b11001001100000;     //407pi/512
   m_cos[407]  =  14'b11011110011100;     //407pi/512
   m_sin[408]  =  14'b11001001101011;     //408pi/512
   m_cos[408]  =  14'b11011110001010;     //408pi/512
   m_sin[409]  =  14'b11001001110111;     //409pi/512
   m_cos[409]  =  14'b11011101111000;     //409pi/512
   m_sin[410]  =  14'b11001010000010;     //410pi/512
   m_cos[410]  =  14'b11011101100110;     //410pi/512
   m_sin[411]  =  14'b11001010001110;     //411pi/512
   m_cos[411]  =  14'b11011101010100;     //411pi/512
   m_sin[412]  =  14'b11001010011001;     //412pi/512
   m_cos[412]  =  14'b11011101000010;     //412pi/512
   m_sin[413]  =  14'b11001010100101;     //413pi/512
   m_cos[413]  =  14'b11011100110000;     //413pi/512
   m_sin[414]  =  14'b11001010110001;     //414pi/512
   m_cos[414]  =  14'b11011100011110;     //414pi/512
   m_sin[415]  =  14'b11001010111101;     //415pi/512
   m_cos[415]  =  14'b11011100001101;     //415pi/512
   m_sin[416]  =  14'b11001011001001;     //416pi/512
   m_cos[416]  =  14'b11011011111011;     //416pi/512
   m_sin[417]  =  14'b11001011010101;     //417pi/512
   m_cos[417]  =  14'b11011011101001;     //417pi/512
   m_sin[418]  =  14'b11001011100001;     //418pi/512
   m_cos[418]  =  14'b11011011011000;     //418pi/512
   m_sin[419]  =  14'b11001011101101;     //419pi/512
   m_cos[419]  =  14'b11011011000110;     //419pi/512
   m_sin[420]  =  14'b11001011111010;     //420pi/512
   m_cos[420]  =  14'b11011010110101;     //420pi/512
   m_sin[421]  =  14'b11001100000110;     //421pi/512
   m_cos[421]  =  14'b11011010100100;     //421pi/512
   m_sin[422]  =  14'b11001100010011;     //422pi/512
   m_cos[422]  =  14'b11011010010010;     //422pi/512
   m_sin[423]  =  14'b11001100011111;     //423pi/512
   m_cos[423]  =  14'b11011010000001;     //423pi/512
   m_sin[424]  =  14'b11001100101100;     //424pi/512
   m_cos[424]  =  14'b11011001110000;     //424pi/512
   m_sin[425]  =  14'b11001100111001;     //425pi/512
   m_cos[425]  =  14'b11011001011111;     //425pi/512
   m_sin[426]  =  14'b11001101000110;     //426pi/512
   m_cos[426]  =  14'b11011001001110;     //426pi/512
   m_sin[427]  =  14'b11001101010011;     //427pi/512
   m_cos[427]  =  14'b11011000111101;     //427pi/512
   m_sin[428]  =  14'b11001101100000;     //428pi/512
   m_cos[428]  =  14'b11011000101100;     //428pi/512
   m_sin[429]  =  14'b11001101101101;     //429pi/512
   m_cos[429]  =  14'b11011000011011;     //429pi/512
   m_sin[430]  =  14'b11001101111010;     //430pi/512
   m_cos[430]  =  14'b11011000001010;     //430pi/512
   m_sin[431]  =  14'b11001110001000;     //431pi/512
   m_cos[431]  =  14'b11010111111010;     //431pi/512
   m_sin[432]  =  14'b11001110010101;     //432pi/512
   m_cos[432]  =  14'b11010111101001;     //432pi/512
   m_sin[433]  =  14'b11001110100011;     //433pi/512
   m_cos[433]  =  14'b11010111011001;     //433pi/512
   m_sin[434]  =  14'b11001110110000;     //434pi/512
   m_cos[434]  =  14'b11010111001000;     //434pi/512
   m_sin[435]  =  14'b11001110111110;     //435pi/512
   m_cos[435]  =  14'b11010110111000;     //435pi/512
   m_sin[436]  =  14'b11001111001100;     //436pi/512
   m_cos[436]  =  14'b11010110100111;     //436pi/512
   m_sin[437]  =  14'b11001111011001;     //437pi/512
   m_cos[437]  =  14'b11010110010111;     //437pi/512
   m_sin[438]  =  14'b11001111100111;     //438pi/512
   m_cos[438]  =  14'b11010110000111;     //438pi/512
   m_sin[439]  =  14'b11001111110101;     //439pi/512
   m_cos[439]  =  14'b11010101110111;     //439pi/512
   m_sin[440]  =  14'b11010000000100;     //440pi/512
   m_cos[440]  =  14'b11010101100111;     //440pi/512
   m_sin[441]  =  14'b11010000010010;     //441pi/512
   m_cos[441]  =  14'b11010101010111;     //441pi/512
   m_sin[442]  =  14'b11010000100000;     //442pi/512
   m_cos[442]  =  14'b11010101000111;     //442pi/512
   m_sin[443]  =  14'b11010000101110;     //443pi/512
   m_cos[443]  =  14'b11010100110111;     //443pi/512
   m_sin[444]  =  14'b11010000111101;     //444pi/512
   m_cos[444]  =  14'b11010100100111;     //444pi/512
   m_sin[445]  =  14'b11010001001011;     //445pi/512
   m_cos[445]  =  14'b11010100011000;     //445pi/512
   m_sin[446]  =  14'b11010001011010;     //446pi/512
   m_cos[446]  =  14'b11010100001000;     //446pi/512
   m_sin[447]  =  14'b11010001101001;     //447pi/512
   m_cos[447]  =  14'b11010011111001;     //447pi/512
   m_sin[448]  =  14'b11010001110111;     //448pi/512
   m_cos[448]  =  14'b11010011101001;     //448pi/512
   m_sin[449]  =  14'b11010010000110;     //449pi/512
   m_cos[449]  =  14'b11010011011010;     //449pi/512
   m_sin[450]  =  14'b11010010010101;     //450pi/512
   m_cos[450]  =  14'b11010011001010;     //450pi/512
   m_sin[451]  =  14'b11010010100100;     //451pi/512
   m_cos[451]  =  14'b11010010111011;     //451pi/512
   m_sin[452]  =  14'b11010010110011;     //452pi/512
   m_cos[452]  =  14'b11010010101100;     //452pi/512
   m_sin[453]  =  14'b11010011000010;     //453pi/512
   m_cos[453]  =  14'b11010010011101;     //453pi/512
   m_sin[454]  =  14'b11010011010010;     //454pi/512
   m_cos[454]  =  14'b11010010001110;     //454pi/512
   m_sin[455]  =  14'b11010011100001;     //455pi/512
   m_cos[455]  =  14'b11010001111111;     //455pi/512
   m_sin[456]  =  14'b11010011110000;     //456pi/512
   m_cos[456]  =  14'b11010001110000;     //456pi/512
   m_sin[457]  =  14'b11010100000000;     //457pi/512
   m_cos[457]  =  14'b11010001100010;     //457pi/512
   m_sin[458]  =  14'b11010100001111;     //458pi/512
   m_cos[458]  =  14'b11010001010011;     //458pi/512
   m_sin[459]  =  14'b11010100011111;     //459pi/512
   m_cos[459]  =  14'b11010001000100;     //459pi/512
   m_sin[460]  =  14'b11010100101111;     //460pi/512
   m_cos[460]  =  14'b11010000110110;     //460pi/512
   m_sin[461]  =  14'b11010100111111;     //461pi/512
   m_cos[461]  =  14'b11010000101000;     //461pi/512
   m_sin[462]  =  14'b11010101001110;     //462pi/512
   m_cos[462]  =  14'b11010000011001;     //462pi/512
   m_sin[463]  =  14'b11010101011110;     //463pi/512
   m_cos[463]  =  14'b11010000001011;     //463pi/512
   m_sin[464]  =  14'b11010101101110;     //464pi/512
   m_cos[464]  =  14'b11001111111101;     //464pi/512
   m_sin[465]  =  14'b11010101111110;     //465pi/512
   m_cos[465]  =  14'b11001111101111;     //465pi/512
   m_sin[466]  =  14'b11010110001111;     //466pi/512
   m_cos[466]  =  14'b11001111100001;     //466pi/512
   m_sin[467]  =  14'b11010110011111;     //467pi/512
   m_cos[467]  =  14'b11001111010011;     //467pi/512
   m_sin[468]  =  14'b11010110101111;     //468pi/512
   m_cos[468]  =  14'b11001111000101;     //468pi/512
   m_sin[469]  =  14'b11010110111111;     //469pi/512
   m_cos[469]  =  14'b11001110110111;     //469pi/512
   m_sin[470]  =  14'b11010111010000;     //470pi/512
   m_cos[470]  =  14'b11001110101010;     //470pi/512
   m_sin[471]  =  14'b11010111100000;     //471pi/512
   m_cos[471]  =  14'b11001110011100;     //471pi/512
   m_sin[472]  =  14'b11010111110001;     //472pi/512
   m_cos[472]  =  14'b11001110001111;     //472pi/512
   m_sin[473]  =  14'b11011000000010;     //473pi/512
   m_cos[473]  =  14'b11001110000001;     //473pi/512
   m_sin[474]  =  14'b11011000010010;     //474pi/512
   m_cos[474]  =  14'b11001101110100;     //474pi/512
   m_sin[475]  =  14'b11011000100011;     //475pi/512
   m_cos[475]  =  14'b11001101100111;     //475pi/512
   m_sin[476]  =  14'b11011000110100;     //476pi/512
   m_cos[476]  =  14'b11001101011010;     //476pi/512
   m_sin[477]  =  14'b11011001000101;     //477pi/512
   m_cos[477]  =  14'b11001101001101;     //477pi/512
   m_sin[478]  =  14'b11011001010110;     //478pi/512
   m_cos[478]  =  14'b11001101000000;     //478pi/512
   m_sin[479]  =  14'b11011001100111;     //479pi/512
   m_cos[479]  =  14'b11001100110011;     //479pi/512
   m_sin[480]  =  14'b11011001111000;     //480pi/512
   m_cos[480]  =  14'b11001100100110;     //480pi/512
   m_sin[481]  =  14'b11011010001001;     //481pi/512
   m_cos[481]  =  14'b11001100011001;     //481pi/512
   m_sin[482]  =  14'b11011010011010;     //482pi/512
   m_cos[482]  =  14'b11001100001101;     //482pi/512
   m_sin[483]  =  14'b11011010101100;     //483pi/512
   m_cos[483]  =  14'b11001100000000;     //483pi/512
   m_sin[484]  =  14'b11011010111101;     //484pi/512
   m_cos[484]  =  14'b11001011110100;     //484pi/512
   m_sin[485]  =  14'b11011011001111;     //485pi/512
   m_cos[485]  =  14'b11001011101000;     //485pi/512
   m_sin[486]  =  14'b11011011100000;     //486pi/512
   m_cos[486]  =  14'b11001011011011;     //486pi/512
   m_sin[487]  =  14'b11011011110010;     //487pi/512
   m_cos[487]  =  14'b11001011001111;     //487pi/512
   m_sin[488]  =  14'b11011100000011;     //488pi/512
   m_cos[488]  =  14'b11001011000011;     //488pi/512
   m_sin[489]  =  14'b11011100010101;     //489pi/512
   m_cos[489]  =  14'b11001010110111;     //489pi/512
   m_sin[490]  =  14'b11011100100111;     //490pi/512
   m_cos[490]  =  14'b11001010101011;     //490pi/512
   m_sin[491]  =  14'b11011100111001;     //491pi/512
   m_cos[491]  =  14'b11001010100000;     //491pi/512
   m_sin[492]  =  14'b11011101001011;     //492pi/512
   m_cos[492]  =  14'b11001010010100;     //492pi/512
   m_sin[493]  =  14'b11011101011101;     //493pi/512
   m_cos[493]  =  14'b11001010001000;     //493pi/512
   m_sin[494]  =  14'b11011101101111;     //494pi/512
   m_cos[494]  =  14'b11001001111101;     //494pi/512
   m_sin[495]  =  14'b11011110000001;     //495pi/512
   m_cos[495]  =  14'b11001001110001;     //495pi/512
   m_sin[496]  =  14'b11011110010011;     //496pi/512
   m_cos[496]  =  14'b11001001100110;     //496pi/512
   m_sin[497]  =  14'b11011110100101;     //497pi/512
   m_cos[497]  =  14'b11001001011011;     //497pi/512
   m_sin[498]  =  14'b11011110110111;     //498pi/512
   m_cos[498]  =  14'b11001001010000;     //498pi/512
   m_sin[499]  =  14'b11011111001001;     //499pi/512
   m_cos[499]  =  14'b11001001000101;     //499pi/512
   m_sin[500]  =  14'b11011111011100;     //500pi/512
   m_cos[500]  =  14'b11001000111010;     //500pi/512
   m_sin[501]  =  14'b11011111101110;     //501pi/512
   m_cos[501]  =  14'b11001000101111;     //501pi/512
   m_sin[502]  =  14'b11100000000001;     //502pi/512
   m_cos[502]  =  14'b11001000100100;     //502pi/512
   m_sin[503]  =  14'b11100000010011;     //503pi/512
   m_cos[503]  =  14'b11001000011010;     //503pi/512
   m_sin[504]  =  14'b11100000100110;     //504pi/512
   m_cos[504]  =  14'b11001000001111;     //504pi/512
   m_sin[505]  =  14'b11100000111000;     //505pi/512
   m_cos[505]  =  14'b11001000000101;     //505pi/512
   m_sin[506]  =  14'b11100001001011;     //506pi/512
   m_cos[506]  =  14'b11000111111010;     //506pi/512
   m_sin[507]  =  14'b11100001011110;     //507pi/512
   m_cos[507]  =  14'b11000111110000;     //507pi/512
   m_sin[508]  =  14'b11100001110001;     //508pi/512
   m_cos[508]  =  14'b11000111100110;     //508pi/512
   m_sin[509]  =  14'b11100010000100;     //509pi/512
   m_cos[509]  =  14'b11000111011100;     //509pi/512
   m_sin[510]  =  14'b11100010010110;     //510pi/512
   m_cos[510]  =  14'b11000111010010;     //510pi/512
   m_sin[511]  =  14'b11100010101001;     //511pi/512
   m_cos[511]  =  14'b11000111001000;     //511pi/512
end

endmodule