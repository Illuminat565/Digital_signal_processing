module  RAM8 #(parameter bit_width=29, N = 16, SIZE = 4)(
    input                              clk,rst_n,
    
    input                              load_data,
    input              [SIZE-1:     0] invert_adr,
    input       signed [bit_width-1:0] Re_i,
    input       signed [bit_width-1:0] Im_i,

    
    input              [SIZE-1:       0]  rd_ptr,
    input                                 en_rd, 

    input              [6:0]             rd_angle_ptr,      

    output reg  signed [bit_width-1:0]  Re_o,
    output reg  signed [bit_width-1:0]  Im_o,
    output reg                          en_radix,
    output  reg signed [13:0]           cos_data,
    output  reg signed [13:0]           sin_data
 );
    reg signed [13:0]  cos  [127:0];
    reg signed [13:0]  sin  [127:0];

    reg  signed  [bit_width-1:0]  mem_Re  [N-1:0];
    reg  signed  [bit_width-1:0]  mem_Im  [N-1:0];

    reg signed [13:0]           cos_temp;
    reg signed [13:0]           sin_temp;

    reg  en_wr_mem;
    reg  en_1;
    reg  en_2;


    


    //------------------------handle read read from MEM----------------------------
        always @(posedge clk) begin
         begin
             if (en_rd) begin
                  Re_o             <= mem_Re[rd_ptr];
                  Im_o             <= mem_Im[rd_ptr];
             end
        end
        end
   //--------------------------handle wirte read from MEM----------------------------
        always @(posedge clk) begin
         begin
           if (load_data)   begin
                  mem_Re[invert_adr] <= Re_i;
                  mem_Im[invert_adr] <= Im_i;    
            end
        end
        end

    //--------------------------------handle reaf tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd ) begin
                  cos_data         <= cos   [rd_angle_ptr];
                  sin_data         <= sin   [rd_angle_ptr];
                  en_radix         <= 1'b1;
             end else en_radix     <= 1'b0;
        end

//-------------------------ROM----------------------------------------------------------
initial begin
   sin[0]  =  14'b00000000000000;     //0pi/128
   cos[0]  =  14'b01000000000000;     //0pi/128
   sin[1]  =  14'b11111110110000;     //1pi/128
   cos[1]  =  14'b00111111111111;     //1pi/128
   sin[2]  =  14'b11111101011111;     //2pi/128
   cos[2]  =  14'b00111111111100;     //2pi/128
   sin[3]  =  14'b11111100001111;     //3pi/128
   cos[3]  =  14'b00111111111000;     //3pi/128
   sin[4]  =  14'b11111010111111;     //4pi/128
   cos[4]  =  14'b00111111110011;     //4pi/128
   sin[5]  =  14'b11111001101111;     //5pi/128
   cos[5]  =  14'b00111111101100;     //5pi/128
   sin[6]  =  14'b11111000011111;     //6pi/128
   cos[6]  =  14'b00111111100011;     //6pi/128
   sin[7]  =  14'b11110111001111;     //7pi/128
   cos[7]  =  14'b00111111011001;     //7pi/128
   sin[8]  =  14'b11110101111111;     //8pi/128
   cos[8]  =  14'b00111111001101;     //8pi/128
   sin[9]  =  14'b11110100110000;     //9pi/128
   cos[9]  =  14'b00111111000000;     //9pi/128
   sin[10]  =  14'b11110011100001;     //10pi/128
   cos[10]  =  14'b00111110110001;     //10pi/128
   sin[11]  =  14'b11110010010010;     //11pi/128
   cos[11]  =  14'b00111110100000;     //11pi/128
   sin[12]  =  14'b11110001000100;     //12pi/128
   cos[12]  =  14'b00111110001110;     //12pi/128
   sin[13]  =  14'b11101111110110;     //13pi/128
   cos[13]  =  14'b00111101111011;     //13pi/128
   sin[14]  =  14'b11101110101000;     //14pi/128
   cos[14]  =  14'b00111101100110;     //14pi/128
   sin[15]  =  14'b11101101011011;     //15pi/128
   cos[15]  =  14'b00111101001111;     //15pi/128
   sin[16]  =  14'b11101100001110;     //16pi/128
   cos[16]  =  14'b00111100110111;     //16pi/128
   sin[17]  =  14'b11101011000010;     //17pi/128
   cos[17]  =  14'b00111100011101;     //17pi/128
   sin[18]  =  14'b11101001110110;     //18pi/128
   cos[18]  =  14'b00111100000010;     //18pi/128
   sin[19]  =  14'b11101000101011;     //19pi/128
   cos[19]  =  14'b00111011100110;     //19pi/128
   sin[20]  =  14'b11100111100001;     //20pi/128
   cos[20]  =  14'b00111011001000;     //20pi/128
   sin[21]  =  14'b11100110010111;     //21pi/128
   cos[21]  =  14'b00111010101000;     //21pi/128
   sin[22]  =  14'b11100101001101;     //22pi/128
   cos[22]  =  14'b00111010000111;     //22pi/128
   sin[23]  =  14'b11100100000100;     //23pi/128
   cos[23]  =  14'b00111001100101;     //23pi/128
   sin[24]  =  14'b11100010111100;     //24pi/128
   cos[24]  =  14'b00111001000001;     //24pi/128
   sin[25]  =  14'b11100001110101;     //25pi/128
   cos[25]  =  14'b00111000011100;     //25pi/128
   sin[26]  =  14'b11100000101111;     //26pi/128
   cos[26]  =  14'b00110111110101;     //26pi/128
   sin[27]  =  14'b11011111101001;     //27pi/128
   cos[27]  =  14'b00110111001101;     //27pi/128
   sin[28]  =  14'b11011110100100;     //28pi/128
   cos[28]  =  14'b00110110100100;     //28pi/128
   sin[29]  =  14'b11011101100000;     //29pi/128
   cos[29]  =  14'b00110101111001;     //29pi/128
   sin[30]  =  14'b11011100011100;     //30pi/128
   cos[30]  =  14'b00110101001101;     //30pi/128
   sin[31]  =  14'b11011011011010;     //31pi/128
   cos[31]  =  14'b00110100100000;     //31pi/128
   sin[32]  =  14'b11011010011000;     //32pi/128
   cos[32]  =  14'b00110011110001;     //32pi/128
   sin[33]  =  14'b11011001011000;     //33pi/128
   cos[33]  =  14'b00110011000001;     //33pi/128
   sin[34]  =  14'b11011000011000;     //34pi/128
   cos[34]  =  14'b00110010010000;     //34pi/128
   sin[35]  =  14'b11010111011010;     //35pi/128
   cos[35]  =  14'b00110001011110;     //35pi/128
   sin[36]  =  14'b11010110011100;     //36pi/128
   cos[36]  =  14'b00110000101010;     //36pi/128
   sin[37]  =  14'b11010101011111;     //37pi/128
   cos[37]  =  14'b00101111110101;     //37pi/128
   sin[38]  =  14'b11010100100100;     //38pi/128
   cos[38]  =  14'b00101110111111;     //38pi/128
   sin[39]  =  14'b11010011101001;     //39pi/128
   cos[39]  =  14'b00101110001000;     //39pi/128
   sin[40]  =  14'b11010010110000;     //40pi/128
   cos[40]  =  14'b00101101010000;     //40pi/128
   sin[41]  =  14'b11010001110111;     //41pi/128
   cos[41]  =  14'b00101100010110;     //41pi/128
   sin[42]  =  14'b11010001000000;     //42pi/128
   cos[42]  =  14'b00101011011100;     //42pi/128
   sin[43]  =  14'b11010000001010;     //43pi/128
   cos[43]  =  14'b00101010100000;     //43pi/128
   sin[44]  =  14'b11001111010101;     //44pi/128
   cos[44]  =  14'b00101001100100;     //44pi/128
   sin[45]  =  14'b11001110100010;     //45pi/128
   cos[45]  =  14'b00101000100110;     //45pi/128
   sin[46]  =  14'b11001101101111;     //46pi/128
   cos[46]  =  14'b00100111100111;     //46pi/128
   sin[47]  =  14'b11001100111110;     //47pi/128
   cos[47]  =  14'b00100110101000;     //47pi/128
   sin[48]  =  14'b11001100001110;     //48pi/128
   cos[48]  =  14'b00100101100111;     //48pi/128
   sin[49]  =  14'b11001011100000;     //49pi/128
   cos[49]  =  14'b00100100100110;     //49pi/128
   sin[50]  =  14'b11001010110010;     //50pi/128
   cos[50]  =  14'b00100011100011;     //50pi/128
   sin[51]  =  14'b11001010000110;     //51pi/128
   cos[51]  =  14'b00100010100000;     //51pi/128
   sin[52]  =  14'b11001001011100;     //52pi/128
   cos[52]  =  14'b00100001011100;     //52pi/128
   sin[53]  =  14'b11001000110010;     //53pi/128
   cos[53]  =  14'b00100000010111;     //53pi/128
   sin[54]  =  14'b11001000001010;     //54pi/128
   cos[54]  =  14'b00011111010001;     //54pi/128
   sin[55]  =  14'b11000111100100;     //55pi/128
   cos[55]  =  14'b00011110001010;     //55pi/128
   sin[56]  =  14'b11000110111110;     //56pi/128
   cos[56]  =  14'b00011101000011;     //56pi/128
   sin[57]  =  14'b11000110011011;     //57pi/128
   cos[57]  =  14'b00011011111011;     //57pi/128
   sin[58]  =  14'b11000101111000;     //58pi/128
   cos[58]  =  14'b00011010110010;     //58pi/128
   sin[59]  =  14'b11000101010111;     //59pi/128
   cos[59]  =  14'b00011001101001;     //59pi/128
   sin[60]  =  14'b11000100111000;     //60pi/128
   cos[60]  =  14'b00011000011111;     //60pi/128
   sin[61]  =  14'b11000100011010;     //61pi/128
   cos[61]  =  14'b00010111010100;     //61pi/128
   sin[62]  =  14'b11000011111101;     //62pi/128
   cos[62]  =  14'b00010110001001;     //62pi/128
   sin[63]  =  14'b11000011100010;     //63pi/128
   cos[63]  =  14'b00010100111101;     //63pi/128
   sin[64]  =  14'b11000011001000;     //64pi/128
   cos[64]  =  14'b00010011110001;     //64pi/128
   sin[65]  =  14'b11000010110000;     //65pi/128
   cos[65]  =  14'b00010010100101;     //65pi/128
   sin[66]  =  14'b11000010011010;     //66pi/128
   cos[66]  =  14'b00010001010111;     //66pi/128
   sin[67]  =  14'b11000010000101;     //67pi/128
   cos[67]  =  14'b00010000001010;     //67pi/128
   sin[68]  =  14'b11000001110001;     //68pi/128
   cos[68]  =  14'b00001110111100;     //68pi/128
   sin[69]  =  14'b11000001011111;     //69pi/128
   cos[69]  =  14'b00001101101101;     //69pi/128
   sin[70]  =  14'b11000001001111;     //70pi/128
   cos[70]  =  14'b00001100011111;     //70pi/128
   sin[71]  =  14'b11000001000000;     //71pi/128
   cos[71]  =  14'b00001011010000;     //71pi/128
   sin[72]  =  14'b11000000110010;     //72pi/128
   cos[72]  =  14'b00001010000000;     //72pi/128
   sin[73]  =  14'b11000000100111;     //73pi/128
   cos[73]  =  14'b00001000110001;     //73pi/128
   sin[74]  =  14'b11000000011100;     //74pi/128
   cos[74]  =  14'b00000111100001;     //74pi/128
   sin[75]  =  14'b11000000010100;     //75pi/128
   cos[75]  =  14'b00000110010001;     //75pi/128
   sin[76]  =  14'b11000000001101;     //76pi/128
   cos[76]  =  14'b00000101000001;     //76pi/128
   sin[77]  =  14'b11000000000111;     //77pi/128
   cos[77]  =  14'b00000011110001;     //77pi/128
   sin[78]  =  14'b11000000000011;     //78pi/128
   cos[78]  =  14'b00000010100000;     //78pi/128
   sin[79]  =  14'b11000000000001;     //79pi/128
   cos[79]  =  14'b00000001010000;     //79pi/128
   sin[80]  =  14'b11000000000000;     //80pi/128
   cos[80]  =  14'b00000000000000;     //80pi/128
   sin[81]  =  14'b11000000000001;     //81pi/128
   cos[81]  =  14'b11111110110000;     //81pi/128
   sin[82]  =  14'b11000000000011;     //82pi/128
   cos[82]  =  14'b11111101011111;     //82pi/128
   sin[83]  =  14'b11000000000111;     //83pi/128
   cos[83]  =  14'b11111100001111;     //83pi/128
   sin[84]  =  14'b11000000001101;     //84pi/128
   cos[84]  =  14'b11111010111111;     //84pi/128
   sin[85]  =  14'b11000000010100;     //85pi/128
   cos[85]  =  14'b11111001101111;     //85pi/128
   sin[86]  =  14'b11000000011100;     //86pi/128
   cos[86]  =  14'b11111000011111;     //86pi/128
   sin[87]  =  14'b11000000100111;     //87pi/128
   cos[87]  =  14'b11110111001111;     //87pi/128
   sin[88]  =  14'b11000000110010;     //88pi/128
   cos[88]  =  14'b11110101111111;     //88pi/128
   sin[89]  =  14'b11000001000000;     //89pi/128
   cos[89]  =  14'b11110100110000;     //89pi/128
   sin[90]  =  14'b11000001001111;     //90pi/128
   cos[90]  =  14'b11110011100001;     //90pi/128
   sin[91]  =  14'b11000001011111;     //91pi/128
   cos[91]  =  14'b11110010010010;     //91pi/128
   sin[92]  =  14'b11000001110001;     //92pi/128
   cos[92]  =  14'b11110001000100;     //92pi/128
   sin[93]  =  14'b11000010000101;     //93pi/128
   cos[93]  =  14'b11101111110110;     //93pi/128
   sin[94]  =  14'b11000010011010;     //94pi/128
   cos[94]  =  14'b11101110101000;     //94pi/128
   sin[95]  =  14'b11000010110000;     //95pi/128
   cos[95]  =  14'b11101101011011;     //95pi/128
   sin[96]  =  14'b11000011001000;     //96pi/128
   cos[96]  =  14'b11101100001110;     //96pi/128
   sin[97]  =  14'b11000011100010;     //97pi/128
   cos[97]  =  14'b11101011000010;     //97pi/128
   sin[98]  =  14'b11000011111101;     //98pi/128
   cos[98]  =  14'b11101001110110;     //98pi/128
   sin[99]  =  14'b11000100011010;     //99pi/128
   cos[99]  =  14'b11101000101011;     //99pi/128
   sin[100]  =  14'b11000100111000;     //100pi/128
   cos[100]  =  14'b11100111100001;     //100pi/128
   sin[101]  =  14'b11000101010111;     //101pi/128
   cos[101]  =  14'b11100110010111;     //101pi/128
   sin[102]  =  14'b11000101111000;     //102pi/128
   cos[102]  =  14'b11100101001101;     //102pi/128
   sin[103]  =  14'b11000110011011;     //103pi/128
   cos[103]  =  14'b11100100000100;     //103pi/128
   sin[104]  =  14'b11000110111110;     //104pi/128
   cos[104]  =  14'b11100010111100;     //104pi/128
   sin[105]  =  14'b11000111100100;     //105pi/128
   cos[105]  =  14'b11100001110101;     //105pi/128
   sin[106]  =  14'b11001000001010;     //106pi/128
   cos[106]  =  14'b11100000101111;     //106pi/128
   sin[107]  =  14'b11001000110010;     //107pi/128
   cos[107]  =  14'b11011111101001;     //107pi/128
   sin[108]  =  14'b11001001011100;     //108pi/128
   cos[108]  =  14'b11011110100100;     //108pi/128
   sin[109]  =  14'b11001010000110;     //109pi/128
   cos[109]  =  14'b11011101100000;     //109pi/128
   sin[110]  =  14'b11001010110010;     //110pi/128
   cos[110]  =  14'b11011100011100;     //110pi/128
   sin[111]  =  14'b11001011100000;     //111pi/128
   cos[111]  =  14'b11011011011010;     //111pi/128
   sin[112]  =  14'b11001100001110;     //112pi/128
   cos[112]  =  14'b11011010011000;     //112pi/128
   sin[113]  =  14'b11001100111110;     //113pi/128
   cos[113]  =  14'b11011001011000;     //113pi/128
   sin[114]  =  14'b11001101101111;     //114pi/128
   cos[114]  =  14'b11011000011000;     //114pi/128
   sin[115]  =  14'b11001110100010;     //115pi/128
   cos[115]  =  14'b11010111011010;     //115pi/128
   sin[116]  =  14'b11001111010101;     //116pi/128
   cos[116]  =  14'b11010110011100;     //116pi/128
   sin[117]  =  14'b11010000001010;     //117pi/128
   cos[117]  =  14'b11010101011111;     //117pi/128
   sin[118]  =  14'b11010001000000;     //118pi/128
   cos[118]  =  14'b11010100100100;     //118pi/128
   sin[119]  =  14'b11010001110111;     //119pi/128
   cos[119]  =  14'b11010011101001;     //119pi/128
   sin[120]  =  14'b11010010110000;     //120pi/128
   cos[120]  =  14'b11010010110000;     //120pi/128
   sin[121]  =  14'b11010011101001;     //121pi/128
   cos[121]  =  14'b11010001110111;     //121pi/128
   sin[122]  =  14'b11010100100100;     //122pi/128
   cos[122]  =  14'b11010001000000;     //122pi/128
   sin[123]  =  14'b11010101011111;     //123pi/128
   cos[123]  =  14'b11010000001010;     //123pi/128
   sin[124]  =  14'b11010110011100;     //124pi/128
   cos[124]  =  14'b11001111010101;     //124pi/128
   sin[125]  =  14'b11010111011010;     //125pi/128
   cos[125]  =  14'b11001110100010;     //125pi/128
   sin[126]  =  14'b11011000011000;     //126pi/128
   cos[126]  =  14'b11001101101111;     //126pi/128
   sin[127]  =  14'b11011001011000;     //127pi/128
   cos[127]  =  14'b11001100111110;     //127pi/128
end

endmodule