module  TWIDLE_14_bit_final_STAGE_2  #(parameter N = 256, SIZE = 8, word_length_tw = 14) (
    input            clk,
    input            en_rd, 
    input   [10:0]   rd_ptr_angle,

    output reg signed [word_length_tw-1:0]   cos_data,
    output reg signed [word_length_tw-1:0]   sin_data
 );

reg signed [word_length_tw-1:0]  cos  [1023:0];
reg signed [word_length_tw-1:0]  sin  [1023:0];



always @(posedge clk) begin
  if (en_rd) begin
    cos_data <= cos [rd_ptr_angle];
    sin_data <= sin [rd_ptr_angle];
  end
end


initial begin
   sin[0]  =  14'b00000000000000;     //0pi/1024
   cos[0]  =  14'b01000000000000;     //0pi/1024
   sin[1]  =  14'b00000000000010;     //0.00019531pi/1024
   cos[1]  =  14'b00111111111111;     //0.00019531pi/1024
   sin[2]  =  14'b00000000000101;     //0.00039063pi/1024
   cos[2]  =  14'b00111111111111;     //0.00039063pi/1024
   sin[3]  =  14'b00000000000111;     //0.00058594pi/1024
   cos[3]  =  14'b00111111111111;     //0.00058594pi/1024
   sin[4]  =  14'b00000000001010;     //0.00078125pi/1024
   cos[4]  =  14'b00111111111111;     //0.00078125pi/1024
   sin[5]  =  14'b00000000001100;     //0.00097656pi/1024
   cos[5]  =  14'b00111111111111;     //0.00097656pi/1024
   sin[6]  =  14'b00000000001111;     //0.0011719pi/1024
   cos[6]  =  14'b00111111111111;     //0.0011719pi/1024
   sin[7]  =  14'b00000000010001;     //0.0013672pi/1024
   cos[7]  =  14'b00111111111111;     //0.0013672pi/1024
   sin[8]  =  14'b00000000010100;     //0.0015625pi/1024
   cos[8]  =  14'b00111111111111;     //0.0015625pi/1024
   sin[9]  =  14'b00000000010110;     //0.0017578pi/1024
   cos[9]  =  14'b00111111111111;     //0.0017578pi/1024
   sin[10]  =  14'b00000000011001;     //0.0019531pi/1024
   cos[10]  =  14'b00111111111111;     //0.0019531pi/1024
   sin[11]  =  14'b00000000011011;     //0.0021484pi/1024
   cos[11]  =  14'b00111111111111;     //0.0021484pi/1024
   sin[12]  =  14'b00000000011110;     //0.0023438pi/1024
   cos[12]  =  14'b00111111111111;     //0.0023438pi/1024
   sin[13]  =  14'b00000000100000;     //0.0025391pi/1024
   cos[13]  =  14'b00111111111111;     //0.0025391pi/1024
   sin[14]  =  14'b00000000100011;     //0.0027344pi/1024
   cos[14]  =  14'b00111111111111;     //0.0027344pi/1024
   sin[15]  =  14'b00000000100101;     //0.0029297pi/1024
   cos[15]  =  14'b00111111111111;     //0.0029297pi/1024
   sin[16]  =  14'b00000000101000;     //0.003125pi/1024
   cos[16]  =  14'b00111111111111;     //0.003125pi/1024
   sin[17]  =  14'b00000000101010;     //0.0033203pi/1024
   cos[17]  =  14'b00111111111111;     //0.0033203pi/1024
   sin[18]  =  14'b00000000101101;     //0.0035156pi/1024
   cos[18]  =  14'b00111111111111;     //0.0035156pi/1024
   sin[19]  =  14'b00000000101111;     //0.0037109pi/1024
   cos[19]  =  14'b00111111111111;     //0.0037109pi/1024
   sin[20]  =  14'b00000000110010;     //0.0039062pi/1024
   cos[20]  =  14'b00111111111111;     //0.0039062pi/1024
   sin[21]  =  14'b00000000110100;     //0.0041016pi/1024
   cos[21]  =  14'b00111111111111;     //0.0041016pi/1024
   sin[22]  =  14'b00000000110111;     //0.0042969pi/1024
   cos[22]  =  14'b00111111111111;     //0.0042969pi/1024
   sin[23]  =  14'b00000000111001;     //0.0044922pi/1024
   cos[23]  =  14'b00111111111111;     //0.0044922pi/1024
   sin[24]  =  14'b00000000111100;     //0.0046875pi/1024
   cos[24]  =  14'b00111111111111;     //0.0046875pi/1024
   sin[25]  =  14'b00000000111110;     //0.0048828pi/1024
   cos[25]  =  14'b00111111111111;     //0.0048828pi/1024
   sin[26]  =  14'b00000001000001;     //0.0050781pi/1024
   cos[26]  =  14'b00111111111111;     //0.0050781pi/1024
   sin[27]  =  14'b00000001000011;     //0.0052734pi/1024
   cos[27]  =  14'b00111111111111;     //0.0052734pi/1024
   sin[28]  =  14'b00000001000110;     //0.0054688pi/1024
   cos[28]  =  14'b00111111111111;     //0.0054688pi/1024
   sin[29]  =  14'b00000001001000;     //0.0056641pi/1024
   cos[29]  =  14'b00111111111111;     //0.0056641pi/1024
   sin[30]  =  14'b00000001001011;     //0.0058594pi/1024
   cos[30]  =  14'b00111111111111;     //0.0058594pi/1024
   sin[31]  =  14'b00000001001101;     //0.0060547pi/1024
   cos[31]  =  14'b00111111111111;     //0.0060547pi/1024
   sin[32]  =  14'b00000001010000;     //0.00625pi/1024
   cos[32]  =  14'b00111111111111;     //0.00625pi/1024
   sin[33]  =  14'b00000001010010;     //0.0064453pi/1024
   cos[33]  =  14'b00111111111111;     //0.0064453pi/1024
   sin[34]  =  14'b00000001010101;     //0.0066406pi/1024
   cos[34]  =  14'b00111111111111;     //0.0066406pi/1024
   sin[35]  =  14'b00000001010111;     //0.0068359pi/1024
   cos[35]  =  14'b00111111111111;     //0.0068359pi/1024
   sin[36]  =  14'b00000001011010;     //0.0070313pi/1024
   cos[36]  =  14'b00111111111111;     //0.0070313pi/1024
   sin[37]  =  14'b00000001011100;     //0.0072266pi/1024
   cos[37]  =  14'b00111111111110;     //0.0072266pi/1024
   sin[38]  =  14'b00000001011111;     //0.0074219pi/1024
   cos[38]  =  14'b00111111111110;     //0.0074219pi/1024
   sin[39]  =  14'b00000001100010;     //0.0076172pi/1024
   cos[39]  =  14'b00111111111110;     //0.0076172pi/1024
   sin[40]  =  14'b00000001100100;     //0.0078125pi/1024
   cos[40]  =  14'b00111111111110;     //0.0078125pi/1024
   sin[41]  =  14'b00000001100111;     //0.0080078pi/1024
   cos[41]  =  14'b00111111111110;     //0.0080078pi/1024
   sin[42]  =  14'b00000001101001;     //0.0082031pi/1024
   cos[42]  =  14'b00111111111110;     //0.0082031pi/1024
   sin[43]  =  14'b00000001101100;     //0.0083984pi/1024
   cos[43]  =  14'b00111111111110;     //0.0083984pi/1024
   sin[44]  =  14'b00000001101110;     //0.0085938pi/1024
   cos[44]  =  14'b00111111111110;     //0.0085938pi/1024
   sin[45]  =  14'b00000001110001;     //0.0087891pi/1024
   cos[45]  =  14'b00111111111110;     //0.0087891pi/1024
   sin[46]  =  14'b00000001110011;     //0.0089844pi/1024
   cos[46]  =  14'b00111111111110;     //0.0089844pi/1024
   sin[47]  =  14'b00000001110110;     //0.0091797pi/1024
   cos[47]  =  14'b00111111111110;     //0.0091797pi/1024
   sin[48]  =  14'b00000001111000;     //0.009375pi/1024
   cos[48]  =  14'b00111111111110;     //0.009375pi/1024
   sin[49]  =  14'b00000001111011;     //0.0095703pi/1024
   cos[49]  =  14'b00111111111110;     //0.0095703pi/1024
   sin[50]  =  14'b00000001111101;     //0.0097656pi/1024
   cos[50]  =  14'b00111111111110;     //0.0097656pi/1024
   sin[51]  =  14'b00000010000000;     //0.0099609pi/1024
   cos[51]  =  14'b00111111111101;     //0.0099609pi/1024
   sin[52]  =  14'b00000010000010;     //0.010156pi/1024
   cos[52]  =  14'b00111111111101;     //0.010156pi/1024
   sin[53]  =  14'b00000010000101;     //0.010352pi/1024
   cos[53]  =  14'b00111111111101;     //0.010352pi/1024
   sin[54]  =  14'b00000010000111;     //0.010547pi/1024
   cos[54]  =  14'b00111111111101;     //0.010547pi/1024
   sin[55]  =  14'b00000010001010;     //0.010742pi/1024
   cos[55]  =  14'b00111111111101;     //0.010742pi/1024
   sin[56]  =  14'b00000010001100;     //0.010938pi/1024
   cos[56]  =  14'b00111111111101;     //0.010938pi/1024
   sin[57]  =  14'b00000010001111;     //0.011133pi/1024
   cos[57]  =  14'b00111111111101;     //0.011133pi/1024
   sin[58]  =  14'b00000010010001;     //0.011328pi/1024
   cos[58]  =  14'b00111111111101;     //0.011328pi/1024
   sin[59]  =  14'b00000010010100;     //0.011523pi/1024
   cos[59]  =  14'b00111111111101;     //0.011523pi/1024
   sin[60]  =  14'b00000010010110;     //0.011719pi/1024
   cos[60]  =  14'b00111111111101;     //0.011719pi/1024
   sin[61]  =  14'b00000010011001;     //0.011914pi/1024
   cos[61]  =  14'b00111111111101;     //0.011914pi/1024
   sin[62]  =  14'b00000010011011;     //0.012109pi/1024
   cos[62]  =  14'b00111111111101;     //0.012109pi/1024
   sin[63]  =  14'b00000010011110;     //0.012305pi/1024
   cos[63]  =  14'b00111111111100;     //0.012305pi/1024
   sin[64]  =  14'b00000010100000;     //0.0125pi/1024
   cos[64]  =  14'b00111111111100;     //0.0125pi/1024
   sin[65]  =  14'b00000010100011;     //0.012695pi/1024
   cos[65]  =  14'b00111111111100;     //0.012695pi/1024
   sin[66]  =  14'b00000010100101;     //0.012891pi/1024
   cos[66]  =  14'b00111111111100;     //0.012891pi/1024
   sin[67]  =  14'b00000010101000;     //0.013086pi/1024
   cos[67]  =  14'b00111111111100;     //0.013086pi/1024
   sin[68]  =  14'b00000010101010;     //0.013281pi/1024
   cos[68]  =  14'b00111111111100;     //0.013281pi/1024
   sin[69]  =  14'b00000010101101;     //0.013477pi/1024
   cos[69]  =  14'b00111111111100;     //0.013477pi/1024
   sin[70]  =  14'b00000010101111;     //0.013672pi/1024
   cos[70]  =  14'b00111111111100;     //0.013672pi/1024
   sin[71]  =  14'b00000010110010;     //0.013867pi/1024
   cos[71]  =  14'b00111111111100;     //0.013867pi/1024
   sin[72]  =  14'b00000010110100;     //0.014063pi/1024
   cos[72]  =  14'b00111111111100;     //0.014063pi/1024
   sin[73]  =  14'b00000010110111;     //0.014258pi/1024
   cos[73]  =  14'b00111111111011;     //0.014258pi/1024
   sin[74]  =  14'b00000010111001;     //0.014453pi/1024
   cos[74]  =  14'b00111111111011;     //0.014453pi/1024
   sin[75]  =  14'b00000010111100;     //0.014648pi/1024
   cos[75]  =  14'b00111111111011;     //0.014648pi/1024
   sin[76]  =  14'b00000010111110;     //0.014844pi/1024
   cos[76]  =  14'b00111111111011;     //0.014844pi/1024
   sin[77]  =  14'b00000011000001;     //0.015039pi/1024
   cos[77]  =  14'b00111111111011;     //0.015039pi/1024
   sin[78]  =  14'b00000011000011;     //0.015234pi/1024
   cos[78]  =  14'b00111111111011;     //0.015234pi/1024
   sin[79]  =  14'b00000011000110;     //0.01543pi/1024
   cos[79]  =  14'b00111111111011;     //0.01543pi/1024
   sin[80]  =  14'b00000011001000;     //0.015625pi/1024
   cos[80]  =  14'b00111111111011;     //0.015625pi/1024
   sin[81]  =  14'b00000011001011;     //0.01582pi/1024
   cos[81]  =  14'b00111111111010;     //0.01582pi/1024
   sin[82]  =  14'b00000011001110;     //0.016016pi/1024
   cos[82]  =  14'b00111111111010;     //0.016016pi/1024
   sin[83]  =  14'b00000011010000;     //0.016211pi/1024
   cos[83]  =  14'b00111111111010;     //0.016211pi/1024
   sin[84]  =  14'b00000011010011;     //0.016406pi/1024
   cos[84]  =  14'b00111111111010;     //0.016406pi/1024
   sin[85]  =  14'b00000011010101;     //0.016602pi/1024
   cos[85]  =  14'b00111111111010;     //0.016602pi/1024
   sin[86]  =  14'b00000011011000;     //0.016797pi/1024
   cos[86]  =  14'b00111111111010;     //0.016797pi/1024
   sin[87]  =  14'b00000011011010;     //0.016992pi/1024
   cos[87]  =  14'b00111111111010;     //0.016992pi/1024
   sin[88]  =  14'b00000011011101;     //0.017188pi/1024
   cos[88]  =  14'b00111111111010;     //0.017188pi/1024
   sin[89]  =  14'b00000011011111;     //0.017383pi/1024
   cos[89]  =  14'b00111111111001;     //0.017383pi/1024
   sin[90]  =  14'b00000011100010;     //0.017578pi/1024
   cos[90]  =  14'b00111111111001;     //0.017578pi/1024
   sin[91]  =  14'b00000011100100;     //0.017773pi/1024
   cos[91]  =  14'b00111111111001;     //0.017773pi/1024
   sin[92]  =  14'b00000011100111;     //0.017969pi/1024
   cos[92]  =  14'b00111111111001;     //0.017969pi/1024
   sin[93]  =  14'b00000011101001;     //0.018164pi/1024
   cos[93]  =  14'b00111111111001;     //0.018164pi/1024
   sin[94]  =  14'b00000011101100;     //0.018359pi/1024
   cos[94]  =  14'b00111111111001;     //0.018359pi/1024
   sin[95]  =  14'b00000011101110;     //0.018555pi/1024
   cos[95]  =  14'b00111111111001;     //0.018555pi/1024
   sin[96]  =  14'b00000011110001;     //0.01875pi/1024
   cos[96]  =  14'b00111111111000;     //0.01875pi/1024
   sin[97]  =  14'b00000011110011;     //0.018945pi/1024
   cos[97]  =  14'b00111111111000;     //0.018945pi/1024
   sin[98]  =  14'b00000011110110;     //0.019141pi/1024
   cos[98]  =  14'b00111111111000;     //0.019141pi/1024
   sin[99]  =  14'b00000011111000;     //0.019336pi/1024
   cos[99]  =  14'b00111111111000;     //0.019336pi/1024
   sin[100]  =  14'b00000011111011;     //0.019531pi/1024
   cos[100]  =  14'b00111111111000;     //0.019531pi/1024
   sin[101]  =  14'b00000011111101;     //0.019727pi/1024
   cos[101]  =  14'b00111111111000;     //0.019727pi/1024
   sin[102]  =  14'b00000100000000;     //0.019922pi/1024
   cos[102]  =  14'b00111111110111;     //0.019922pi/1024
   sin[103]  =  14'b00000100000010;     //0.020117pi/1024
   cos[103]  =  14'b00111111110111;     //0.020117pi/1024
   sin[104]  =  14'b00000100000101;     //0.020313pi/1024
   cos[104]  =  14'b00111111110111;     //0.020313pi/1024
   sin[105]  =  14'b00000100000111;     //0.020508pi/1024
   cos[105]  =  14'b00111111110111;     //0.020508pi/1024
   sin[106]  =  14'b00000100001010;     //0.020703pi/1024
   cos[106]  =  14'b00111111110111;     //0.020703pi/1024
   sin[107]  =  14'b00000100001100;     //0.020898pi/1024
   cos[107]  =  14'b00111111110111;     //0.020898pi/1024
   sin[108]  =  14'b00000100001111;     //0.021094pi/1024
   cos[108]  =  14'b00111111110111;     //0.021094pi/1024
   sin[109]  =  14'b00000100010001;     //0.021289pi/1024
   cos[109]  =  14'b00111111110110;     //0.021289pi/1024
   sin[110]  =  14'b00000100010100;     //0.021484pi/1024
   cos[110]  =  14'b00111111110110;     //0.021484pi/1024
   sin[111]  =  14'b00000100010110;     //0.02168pi/1024
   cos[111]  =  14'b00111111110110;     //0.02168pi/1024
   sin[112]  =  14'b00000100011001;     //0.021875pi/1024
   cos[112]  =  14'b00111111110110;     //0.021875pi/1024
   sin[113]  =  14'b00000100011011;     //0.02207pi/1024
   cos[113]  =  14'b00111111110110;     //0.02207pi/1024
   sin[114]  =  14'b00000100011110;     //0.022266pi/1024
   cos[114]  =  14'b00111111110101;     //0.022266pi/1024
   sin[115]  =  14'b00000100100000;     //0.022461pi/1024
   cos[115]  =  14'b00111111110101;     //0.022461pi/1024
   sin[116]  =  14'b00000100100011;     //0.022656pi/1024
   cos[116]  =  14'b00111111110101;     //0.022656pi/1024
   sin[117]  =  14'b00000100100101;     //0.022852pi/1024
   cos[117]  =  14'b00111111110101;     //0.022852pi/1024
   sin[118]  =  14'b00000100101000;     //0.023047pi/1024
   cos[118]  =  14'b00111111110101;     //0.023047pi/1024
   sin[119]  =  14'b00000100101010;     //0.023242pi/1024
   cos[119]  =  14'b00111111110101;     //0.023242pi/1024
   sin[120]  =  14'b00000100101101;     //0.023438pi/1024
   cos[120]  =  14'b00111111110100;     //0.023438pi/1024
   sin[121]  =  14'b00000100101111;     //0.023633pi/1024
   cos[121]  =  14'b00111111110100;     //0.023633pi/1024
   sin[122]  =  14'b00000100110010;     //0.023828pi/1024
   cos[122]  =  14'b00111111110100;     //0.023828pi/1024
   sin[123]  =  14'b00000100110100;     //0.024023pi/1024
   cos[123]  =  14'b00111111110100;     //0.024023pi/1024
   sin[124]  =  14'b00000100110111;     //0.024219pi/1024
   cos[124]  =  14'b00111111110100;     //0.024219pi/1024
   sin[125]  =  14'b00000100111001;     //0.024414pi/1024
   cos[125]  =  14'b00111111110011;     //0.024414pi/1024
   sin[126]  =  14'b00000100111100;     //0.024609pi/1024
   cos[126]  =  14'b00111111110011;     //0.024609pi/1024
   sin[127]  =  14'b00000100111110;     //0.024805pi/1024
   cos[127]  =  14'b00111111110011;     //0.024805pi/1024
   sin[128]  =  14'b00000101000001;     //0.025pi/1024
   cos[128]  =  14'b00111111110011;     //0.025pi/1024
   sin[129]  =  14'b00000101000011;     //0.025195pi/1024
   cos[129]  =  14'b00111111110011;     //0.025195pi/1024
   sin[130]  =  14'b00000101000110;     //0.025391pi/1024
   cos[130]  =  14'b00111111110010;     //0.025391pi/1024
   sin[131]  =  14'b00000101001000;     //0.025586pi/1024
   cos[131]  =  14'b00111111110010;     //0.025586pi/1024
   sin[132]  =  14'b00000101001011;     //0.025781pi/1024
   cos[132]  =  14'b00111111110010;     //0.025781pi/1024
   sin[133]  =  14'b00000101001101;     //0.025977pi/1024
   cos[133]  =  14'b00111111110010;     //0.025977pi/1024
   sin[134]  =  14'b00000101010000;     //0.026172pi/1024
   cos[134]  =  14'b00111111110010;     //0.026172pi/1024
   sin[135]  =  14'b00000101010010;     //0.026367pi/1024
   cos[135]  =  14'b00111111110001;     //0.026367pi/1024
   sin[136]  =  14'b00000101010101;     //0.026563pi/1024
   cos[136]  =  14'b00111111110001;     //0.026563pi/1024
   sin[137]  =  14'b00000101010111;     //0.026758pi/1024
   cos[137]  =  14'b00111111110001;     //0.026758pi/1024
   sin[138]  =  14'b00000101011010;     //0.026953pi/1024
   cos[138]  =  14'b00111111110001;     //0.026953pi/1024
   sin[139]  =  14'b00000101011100;     //0.027148pi/1024
   cos[139]  =  14'b00111111110001;     //0.027148pi/1024
   sin[140]  =  14'b00000101011111;     //0.027344pi/1024
   cos[140]  =  14'b00111111110000;     //0.027344pi/1024
   sin[141]  =  14'b00000101100001;     //0.027539pi/1024
   cos[141]  =  14'b00111111110000;     //0.027539pi/1024
   sin[142]  =  14'b00000101100100;     //0.027734pi/1024
   cos[142]  =  14'b00111111110000;     //0.027734pi/1024
   sin[143]  =  14'b00000101100110;     //0.02793pi/1024
   cos[143]  =  14'b00111111110000;     //0.02793pi/1024
   sin[144]  =  14'b00000101101001;     //0.028125pi/1024
   cos[144]  =  14'b00111111110000;     //0.028125pi/1024
   sin[145]  =  14'b00000101101011;     //0.02832pi/1024
   cos[145]  =  14'b00111111101111;     //0.02832pi/1024
   sin[146]  =  14'b00000101101110;     //0.028516pi/1024
   cos[146]  =  14'b00111111101111;     //0.028516pi/1024
   sin[147]  =  14'b00000101110000;     //0.028711pi/1024
   cos[147]  =  14'b00111111101111;     //0.028711pi/1024
   sin[148]  =  14'b00000101110011;     //0.028906pi/1024
   cos[148]  =  14'b00111111101111;     //0.028906pi/1024
   sin[149]  =  14'b00000101110101;     //0.029102pi/1024
   cos[149]  =  14'b00111111101110;     //0.029102pi/1024
   sin[150]  =  14'b00000101111000;     //0.029297pi/1024
   cos[150]  =  14'b00111111101110;     //0.029297pi/1024
   sin[151]  =  14'b00000101111010;     //0.029492pi/1024
   cos[151]  =  14'b00111111101110;     //0.029492pi/1024
   sin[152]  =  14'b00000101111101;     //0.029688pi/1024
   cos[152]  =  14'b00111111101110;     //0.029688pi/1024
   sin[153]  =  14'b00000101111111;     //0.029883pi/1024
   cos[153]  =  14'b00111111101101;     //0.029883pi/1024
   sin[154]  =  14'b00000110000010;     //0.030078pi/1024
   cos[154]  =  14'b00111111101101;     //0.030078pi/1024
   sin[155]  =  14'b00000110000100;     //0.030273pi/1024
   cos[155]  =  14'b00111111101101;     //0.030273pi/1024
   sin[156]  =  14'b00000110000111;     //0.030469pi/1024
   cos[156]  =  14'b00111111101101;     //0.030469pi/1024
   sin[157]  =  14'b00000110001001;     //0.030664pi/1024
   cos[157]  =  14'b00111111101101;     //0.030664pi/1024
   sin[158]  =  14'b00000110001100;     //0.030859pi/1024
   cos[158]  =  14'b00111111101100;     //0.030859pi/1024
   sin[159]  =  14'b00000110001110;     //0.031055pi/1024
   cos[159]  =  14'b00111111101100;     //0.031055pi/1024
   sin[160]  =  14'b00000110010001;     //0.03125pi/1024
   cos[160]  =  14'b00111111101100;     //0.03125pi/1024
   sin[161]  =  14'b00000110010011;     //0.031445pi/1024
   cos[161]  =  14'b00111111101100;     //0.031445pi/1024
   sin[162]  =  14'b00000110010110;     //0.031641pi/1024
   cos[162]  =  14'b00111111101011;     //0.031641pi/1024
   sin[163]  =  14'b00000110011000;     //0.031836pi/1024
   cos[163]  =  14'b00111111101011;     //0.031836pi/1024
   sin[164]  =  14'b00000110011011;     //0.032031pi/1024
   cos[164]  =  14'b00111111101011;     //0.032031pi/1024
   sin[165]  =  14'b00000110011101;     //0.032227pi/1024
   cos[165]  =  14'b00111111101011;     //0.032227pi/1024
   sin[166]  =  14'b00000110100000;     //0.032422pi/1024
   cos[166]  =  14'b00111111101010;     //0.032422pi/1024
   sin[167]  =  14'b00000110100010;     //0.032617pi/1024
   cos[167]  =  14'b00111111101010;     //0.032617pi/1024
   sin[168]  =  14'b00000110100101;     //0.032813pi/1024
   cos[168]  =  14'b00111111101010;     //0.032813pi/1024
   sin[169]  =  14'b00000110100111;     //0.033008pi/1024
   cos[169]  =  14'b00111111101001;     //0.033008pi/1024
   sin[170]  =  14'b00000110101010;     //0.033203pi/1024
   cos[170]  =  14'b00111111101001;     //0.033203pi/1024
   sin[171]  =  14'b00000110101100;     //0.033398pi/1024
   cos[171]  =  14'b00111111101001;     //0.033398pi/1024
   sin[172]  =  14'b00000110101111;     //0.033594pi/1024
   cos[172]  =  14'b00111111101001;     //0.033594pi/1024
   sin[173]  =  14'b00000110110001;     //0.033789pi/1024
   cos[173]  =  14'b00111111101000;     //0.033789pi/1024
   sin[174]  =  14'b00000110110100;     //0.033984pi/1024
   cos[174]  =  14'b00111111101000;     //0.033984pi/1024
   sin[175]  =  14'b00000110110110;     //0.03418pi/1024
   cos[175]  =  14'b00111111101000;     //0.03418pi/1024
   sin[176]  =  14'b00000110111001;     //0.034375pi/1024
   cos[176]  =  14'b00111111101000;     //0.034375pi/1024
   sin[177]  =  14'b00000110111011;     //0.03457pi/1024
   cos[177]  =  14'b00111111100111;     //0.03457pi/1024
   sin[178]  =  14'b00000110111110;     //0.034766pi/1024
   cos[178]  =  14'b00111111100111;     //0.034766pi/1024
   sin[179]  =  14'b00000111000000;     //0.034961pi/1024
   cos[179]  =  14'b00111111100111;     //0.034961pi/1024
   sin[180]  =  14'b00000111000011;     //0.035156pi/1024
   cos[180]  =  14'b00111111100111;     //0.035156pi/1024
   sin[181]  =  14'b00000111000101;     //0.035352pi/1024
   cos[181]  =  14'b00111111100110;     //0.035352pi/1024
   sin[182]  =  14'b00000111001000;     //0.035547pi/1024
   cos[182]  =  14'b00111111100110;     //0.035547pi/1024
   sin[183]  =  14'b00000111001010;     //0.035742pi/1024
   cos[183]  =  14'b00111111100110;     //0.035742pi/1024
   sin[184]  =  14'b00000111001101;     //0.035938pi/1024
   cos[184]  =  14'b00111111100101;     //0.035938pi/1024
   sin[185]  =  14'b00000111001111;     //0.036133pi/1024
   cos[185]  =  14'b00111111100101;     //0.036133pi/1024
   sin[186]  =  14'b00000111010010;     //0.036328pi/1024
   cos[186]  =  14'b00111111100101;     //0.036328pi/1024
   sin[187]  =  14'b00000111010100;     //0.036523pi/1024
   cos[187]  =  14'b00111111100101;     //0.036523pi/1024
   sin[188]  =  14'b00000111010111;     //0.036719pi/1024
   cos[188]  =  14'b00111111100100;     //0.036719pi/1024
   sin[189]  =  14'b00000111011001;     //0.036914pi/1024
   cos[189]  =  14'b00111111100100;     //0.036914pi/1024
   sin[190]  =  14'b00000111011100;     //0.037109pi/1024
   cos[190]  =  14'b00111111100100;     //0.037109pi/1024
   sin[191]  =  14'b00000111011110;     //0.037305pi/1024
   cos[191]  =  14'b00111111100011;     //0.037305pi/1024
   sin[192]  =  14'b00000111100001;     //0.0375pi/1024
   cos[192]  =  14'b00111111100011;     //0.0375pi/1024
   sin[193]  =  14'b00000111100011;     //0.037695pi/1024
   cos[193]  =  14'b00111111100011;     //0.037695pi/1024
   sin[194]  =  14'b00000111100110;     //0.037891pi/1024
   cos[194]  =  14'b00111111100011;     //0.037891pi/1024
   sin[195]  =  14'b00000111101000;     //0.038086pi/1024
   cos[195]  =  14'b00111111100010;     //0.038086pi/1024
   sin[196]  =  14'b00000111101011;     //0.038281pi/1024
   cos[196]  =  14'b00111111100010;     //0.038281pi/1024
   sin[197]  =  14'b00000111101101;     //0.038477pi/1024
   cos[197]  =  14'b00111111100010;     //0.038477pi/1024
   sin[198]  =  14'b00000111110000;     //0.038672pi/1024
   cos[198]  =  14'b00111111100001;     //0.038672pi/1024
   sin[199]  =  14'b00000111110010;     //0.038867pi/1024
   cos[199]  =  14'b00111111100001;     //0.038867pi/1024
   sin[200]  =  14'b00000111110101;     //0.039062pi/1024
   cos[200]  =  14'b00111111100001;     //0.039062pi/1024
   sin[201]  =  14'b00000111110111;     //0.039258pi/1024
   cos[201]  =  14'b00111111100000;     //0.039258pi/1024
   sin[202]  =  14'b00000111111010;     //0.039453pi/1024
   cos[202]  =  14'b00111111100000;     //0.039453pi/1024
   sin[203]  =  14'b00000111111100;     //0.039648pi/1024
   cos[203]  =  14'b00111111100000;     //0.039648pi/1024
   sin[204]  =  14'b00000111111111;     //0.039844pi/1024
   cos[204]  =  14'b00111111011111;     //0.039844pi/1024
   sin[205]  =  14'b00001000000001;     //0.040039pi/1024
   cos[205]  =  14'b00111111011111;     //0.040039pi/1024
   sin[206]  =  14'b00001000000100;     //0.040234pi/1024
   cos[206]  =  14'b00111111011111;     //0.040234pi/1024
   sin[207]  =  14'b00001000000110;     //0.04043pi/1024
   cos[207]  =  14'b00111111011111;     //0.04043pi/1024
   sin[208]  =  14'b00001000001001;     //0.040625pi/1024
   cos[208]  =  14'b00111111011110;     //0.040625pi/1024
   sin[209]  =  14'b00001000001011;     //0.04082pi/1024
   cos[209]  =  14'b00111111011110;     //0.04082pi/1024
   sin[210]  =  14'b00001000001110;     //0.041016pi/1024
   cos[210]  =  14'b00111111011110;     //0.041016pi/1024
   sin[211]  =  14'b00001000010000;     //0.041211pi/1024
   cos[211]  =  14'b00111111011101;     //0.041211pi/1024
   sin[212]  =  14'b00001000010011;     //0.041406pi/1024
   cos[212]  =  14'b00111111011101;     //0.041406pi/1024
   sin[213]  =  14'b00001000010101;     //0.041602pi/1024
   cos[213]  =  14'b00111111011101;     //0.041602pi/1024
   sin[214]  =  14'b00001000011000;     //0.041797pi/1024
   cos[214]  =  14'b00111111011100;     //0.041797pi/1024
   sin[215]  =  14'b00001000011010;     //0.041992pi/1024
   cos[215]  =  14'b00111111011100;     //0.041992pi/1024
   sin[216]  =  14'b00001000011101;     //0.042188pi/1024
   cos[216]  =  14'b00111111011100;     //0.042188pi/1024
   sin[217]  =  14'b00001000011111;     //0.042383pi/1024
   cos[217]  =  14'b00111111011011;     //0.042383pi/1024
   sin[218]  =  14'b00001000100010;     //0.042578pi/1024
   cos[218]  =  14'b00111111011011;     //0.042578pi/1024
   sin[219]  =  14'b00001000100100;     //0.042773pi/1024
   cos[219]  =  14'b00111111011011;     //0.042773pi/1024
   sin[220]  =  14'b00001000100111;     //0.042969pi/1024
   cos[220]  =  14'b00111111011010;     //0.042969pi/1024
   sin[221]  =  14'b00001000101001;     //0.043164pi/1024
   cos[221]  =  14'b00111111011010;     //0.043164pi/1024
   sin[222]  =  14'b00001000101100;     //0.043359pi/1024
   cos[222]  =  14'b00111111011010;     //0.043359pi/1024
   sin[223]  =  14'b00001000101110;     //0.043555pi/1024
   cos[223]  =  14'b00111111011001;     //0.043555pi/1024
   sin[224]  =  14'b00001000110001;     //0.04375pi/1024
   cos[224]  =  14'b00111111011001;     //0.04375pi/1024
   sin[225]  =  14'b00001000110011;     //0.043945pi/1024
   cos[225]  =  14'b00111111011001;     //0.043945pi/1024
   sin[226]  =  14'b00001000110110;     //0.044141pi/1024
   cos[226]  =  14'b00111111011000;     //0.044141pi/1024
   sin[227]  =  14'b00001000111000;     //0.044336pi/1024
   cos[227]  =  14'b00111111011000;     //0.044336pi/1024
   sin[228]  =  14'b00001000111011;     //0.044531pi/1024
   cos[228]  =  14'b00111111010111;     //0.044531pi/1024
   sin[229]  =  14'b00001000111101;     //0.044727pi/1024
   cos[229]  =  14'b00111111010111;     //0.044727pi/1024
   sin[230]  =  14'b00001001000000;     //0.044922pi/1024
   cos[230]  =  14'b00111111010111;     //0.044922pi/1024
   sin[231]  =  14'b00001001000010;     //0.045117pi/1024
   cos[231]  =  14'b00111111010110;     //0.045117pi/1024
   sin[232]  =  14'b00001001000101;     //0.045313pi/1024
   cos[232]  =  14'b00111111010110;     //0.045313pi/1024
   sin[233]  =  14'b00001001000111;     //0.045508pi/1024
   cos[233]  =  14'b00111111010110;     //0.045508pi/1024
   sin[234]  =  14'b00001001001010;     //0.045703pi/1024
   cos[234]  =  14'b00111111010101;     //0.045703pi/1024
   sin[235]  =  14'b00001001001100;     //0.045898pi/1024
   cos[235]  =  14'b00111111010101;     //0.045898pi/1024
   sin[236]  =  14'b00001001001111;     //0.046094pi/1024
   cos[236]  =  14'b00111111010101;     //0.046094pi/1024
   sin[237]  =  14'b00001001010001;     //0.046289pi/1024
   cos[237]  =  14'b00111111010100;     //0.046289pi/1024
   sin[238]  =  14'b00001001010100;     //0.046484pi/1024
   cos[238]  =  14'b00111111010100;     //0.046484pi/1024
   sin[239]  =  14'b00001001010110;     //0.04668pi/1024
   cos[239]  =  14'b00111111010100;     //0.04668pi/1024
   sin[240]  =  14'b00001001011001;     //0.046875pi/1024
   cos[240]  =  14'b00111111010011;     //0.046875pi/1024
   sin[241]  =  14'b00001001011011;     //0.04707pi/1024
   cos[241]  =  14'b00111111010011;     //0.04707pi/1024
   sin[242]  =  14'b00001001011101;     //0.047266pi/1024
   cos[242]  =  14'b00111111010010;     //0.047266pi/1024
   sin[243]  =  14'b00001001100000;     //0.047461pi/1024
   cos[243]  =  14'b00111111010010;     //0.047461pi/1024
   sin[244]  =  14'b00001001100010;     //0.047656pi/1024
   cos[244]  =  14'b00111111010010;     //0.047656pi/1024
   sin[245]  =  14'b00001001100101;     //0.047852pi/1024
   cos[245]  =  14'b00111111010001;     //0.047852pi/1024
   sin[246]  =  14'b00001001100111;     //0.048047pi/1024
   cos[246]  =  14'b00111111010001;     //0.048047pi/1024
   sin[247]  =  14'b00001001101010;     //0.048242pi/1024
   cos[247]  =  14'b00111111010001;     //0.048242pi/1024
   sin[248]  =  14'b00001001101100;     //0.048438pi/1024
   cos[248]  =  14'b00111111010000;     //0.048438pi/1024
   sin[249]  =  14'b00001001101111;     //0.048633pi/1024
   cos[249]  =  14'b00111111010000;     //0.048633pi/1024
   sin[250]  =  14'b00001001110001;     //0.048828pi/1024
   cos[250]  =  14'b00111111001111;     //0.048828pi/1024
   sin[251]  =  14'b00001001110100;     //0.049023pi/1024
   cos[251]  =  14'b00111111001111;     //0.049023pi/1024
   sin[252]  =  14'b00001001110110;     //0.049219pi/1024
   cos[252]  =  14'b00111111001111;     //0.049219pi/1024
   sin[253]  =  14'b00001001111001;     //0.049414pi/1024
   cos[253]  =  14'b00111111001110;     //0.049414pi/1024
   sin[254]  =  14'b00001001111011;     //0.049609pi/1024
   cos[254]  =  14'b00111111001110;     //0.049609pi/1024
   sin[255]  =  14'b00001001111110;     //0.049805pi/1024
   cos[255]  =  14'b00111111001101;     //0.049805pi/1024
   sin[256]  =  14'b00001010000000;     //0.05pi/1024
   cos[256]  =  14'b00111111001101;     //0.05pi/1024
   sin[257]  =  14'b00001010000011;     //0.050195pi/1024
   cos[257]  =  14'b00111111001101;     //0.050195pi/1024
   sin[258]  =  14'b00001010000101;     //0.050391pi/1024
   cos[258]  =  14'b00111111001100;     //0.050391pi/1024
   sin[259]  =  14'b00001010001000;     //0.050586pi/1024
   cos[259]  =  14'b00111111001100;     //0.050586pi/1024
   sin[260]  =  14'b00001010001010;     //0.050781pi/1024
   cos[260]  =  14'b00111111001011;     //0.050781pi/1024
   sin[261]  =  14'b00001010001101;     //0.050977pi/1024
   cos[261]  =  14'b00111111001011;     //0.050977pi/1024
   sin[262]  =  14'b00001010001111;     //0.051172pi/1024
   cos[262]  =  14'b00111111001011;     //0.051172pi/1024
   sin[263]  =  14'b00001010010010;     //0.051367pi/1024
   cos[263]  =  14'b00111111001010;     //0.051367pi/1024
   sin[264]  =  14'b00001010010100;     //0.051563pi/1024
   cos[264]  =  14'b00111111001010;     //0.051563pi/1024
   sin[265]  =  14'b00001010010111;     //0.051758pi/1024
   cos[265]  =  14'b00111111001001;     //0.051758pi/1024
   sin[266]  =  14'b00001010011001;     //0.051953pi/1024
   cos[266]  =  14'b00111111001001;     //0.051953pi/1024
   sin[267]  =  14'b00001010011100;     //0.052148pi/1024
   cos[267]  =  14'b00111111001001;     //0.052148pi/1024
   sin[268]  =  14'b00001010011110;     //0.052344pi/1024
   cos[268]  =  14'b00111111001000;     //0.052344pi/1024
   sin[269]  =  14'b00001010100001;     //0.052539pi/1024
   cos[269]  =  14'b00111111001000;     //0.052539pi/1024
   sin[270]  =  14'b00001010100011;     //0.052734pi/1024
   cos[270]  =  14'b00111111000111;     //0.052734pi/1024
   sin[271]  =  14'b00001010100101;     //0.05293pi/1024
   cos[271]  =  14'b00111111000111;     //0.05293pi/1024
   sin[272]  =  14'b00001010101000;     //0.053125pi/1024
   cos[272]  =  14'b00111111000111;     //0.053125pi/1024
   sin[273]  =  14'b00001010101010;     //0.05332pi/1024
   cos[273]  =  14'b00111111000110;     //0.05332pi/1024
   sin[274]  =  14'b00001010101101;     //0.053516pi/1024
   cos[274]  =  14'b00111111000110;     //0.053516pi/1024
   sin[275]  =  14'b00001010101111;     //0.053711pi/1024
   cos[275]  =  14'b00111111000101;     //0.053711pi/1024
   sin[276]  =  14'b00001010110010;     //0.053906pi/1024
   cos[276]  =  14'b00111111000101;     //0.053906pi/1024
   sin[277]  =  14'b00001010110100;     //0.054102pi/1024
   cos[277]  =  14'b00111111000100;     //0.054102pi/1024
   sin[278]  =  14'b00001010110111;     //0.054297pi/1024
   cos[278]  =  14'b00111111000100;     //0.054297pi/1024
   sin[279]  =  14'b00001010111001;     //0.054492pi/1024
   cos[279]  =  14'b00111111000100;     //0.054492pi/1024
   sin[280]  =  14'b00001010111100;     //0.054688pi/1024
   cos[280]  =  14'b00111111000011;     //0.054688pi/1024
   sin[281]  =  14'b00001010111110;     //0.054883pi/1024
   cos[281]  =  14'b00111111000011;     //0.054883pi/1024
   sin[282]  =  14'b00001011000001;     //0.055078pi/1024
   cos[282]  =  14'b00111111000010;     //0.055078pi/1024
   sin[283]  =  14'b00001011000011;     //0.055273pi/1024
   cos[283]  =  14'b00111111000010;     //0.055273pi/1024
   sin[284]  =  14'b00001011000110;     //0.055469pi/1024
   cos[284]  =  14'b00111111000001;     //0.055469pi/1024
   sin[285]  =  14'b00001011001000;     //0.055664pi/1024
   cos[285]  =  14'b00111111000001;     //0.055664pi/1024
   sin[286]  =  14'b00001011001011;     //0.055859pi/1024
   cos[286]  =  14'b00111111000001;     //0.055859pi/1024
   sin[287]  =  14'b00001011001101;     //0.056055pi/1024
   cos[287]  =  14'b00111111000000;     //0.056055pi/1024
   sin[288]  =  14'b00001011010000;     //0.05625pi/1024
   cos[288]  =  14'b00111111000000;     //0.05625pi/1024
   sin[289]  =  14'b00001011010010;     //0.056445pi/1024
   cos[289]  =  14'b00111110111111;     //0.056445pi/1024
   sin[290]  =  14'b00001011010101;     //0.056641pi/1024
   cos[290]  =  14'b00111110111111;     //0.056641pi/1024
   sin[291]  =  14'b00001011010111;     //0.056836pi/1024
   cos[291]  =  14'b00111110111110;     //0.056836pi/1024
   sin[292]  =  14'b00001011011001;     //0.057031pi/1024
   cos[292]  =  14'b00111110111110;     //0.057031pi/1024
   sin[293]  =  14'b00001011011100;     //0.057227pi/1024
   cos[293]  =  14'b00111110111101;     //0.057227pi/1024
   sin[294]  =  14'b00001011011110;     //0.057422pi/1024
   cos[294]  =  14'b00111110111101;     //0.057422pi/1024
   sin[295]  =  14'b00001011100001;     //0.057617pi/1024
   cos[295]  =  14'b00111110111101;     //0.057617pi/1024
   sin[296]  =  14'b00001011100011;     //0.057813pi/1024
   cos[296]  =  14'b00111110111100;     //0.057813pi/1024
   sin[297]  =  14'b00001011100110;     //0.058008pi/1024
   cos[297]  =  14'b00111110111100;     //0.058008pi/1024
   sin[298]  =  14'b00001011101000;     //0.058203pi/1024
   cos[298]  =  14'b00111110111011;     //0.058203pi/1024
   sin[299]  =  14'b00001011101011;     //0.058398pi/1024
   cos[299]  =  14'b00111110111011;     //0.058398pi/1024
   sin[300]  =  14'b00001011101101;     //0.058594pi/1024
   cos[300]  =  14'b00111110111010;     //0.058594pi/1024
   sin[301]  =  14'b00001011110000;     //0.058789pi/1024
   cos[301]  =  14'b00111110111010;     //0.058789pi/1024
   sin[302]  =  14'b00001011110010;     //0.058984pi/1024
   cos[302]  =  14'b00111110111001;     //0.058984pi/1024
   sin[303]  =  14'b00001011110101;     //0.05918pi/1024
   cos[303]  =  14'b00111110111001;     //0.05918pi/1024
   sin[304]  =  14'b00001011110111;     //0.059375pi/1024
   cos[304]  =  14'b00111110111000;     //0.059375pi/1024
   sin[305]  =  14'b00001011111010;     //0.05957pi/1024
   cos[305]  =  14'b00111110111000;     //0.05957pi/1024
   sin[306]  =  14'b00001011111100;     //0.059766pi/1024
   cos[306]  =  14'b00111110111000;     //0.059766pi/1024
   sin[307]  =  14'b00001011111111;     //0.059961pi/1024
   cos[307]  =  14'b00111110110111;     //0.059961pi/1024
   sin[308]  =  14'b00001100000001;     //0.060156pi/1024
   cos[308]  =  14'b00111110110111;     //0.060156pi/1024
   sin[309]  =  14'b00001100000011;     //0.060352pi/1024
   cos[309]  =  14'b00111110110110;     //0.060352pi/1024
   sin[310]  =  14'b00001100000110;     //0.060547pi/1024
   cos[310]  =  14'b00111110110110;     //0.060547pi/1024
   sin[311]  =  14'b00001100001000;     //0.060742pi/1024
   cos[311]  =  14'b00111110110101;     //0.060742pi/1024
   sin[312]  =  14'b00001100001011;     //0.060938pi/1024
   cos[312]  =  14'b00111110110101;     //0.060938pi/1024
   sin[313]  =  14'b00001100001101;     //0.061133pi/1024
   cos[313]  =  14'b00111110110100;     //0.061133pi/1024
   sin[314]  =  14'b00001100010000;     //0.061328pi/1024
   cos[314]  =  14'b00111110110100;     //0.061328pi/1024
   sin[315]  =  14'b00001100010010;     //0.061523pi/1024
   cos[315]  =  14'b00111110110011;     //0.061523pi/1024
   sin[316]  =  14'b00001100010101;     //0.061719pi/1024
   cos[316]  =  14'b00111110110011;     //0.061719pi/1024
   sin[317]  =  14'b00001100010111;     //0.061914pi/1024
   cos[317]  =  14'b00111110110010;     //0.061914pi/1024
   sin[318]  =  14'b00001100011010;     //0.062109pi/1024
   cos[318]  =  14'b00111110110010;     //0.062109pi/1024
   sin[319]  =  14'b00001100011100;     //0.062305pi/1024
   cos[319]  =  14'b00111110110001;     //0.062305pi/1024
   sin[320]  =  14'b00001100011111;     //0.0625pi/1024
   cos[320]  =  14'b00111110110001;     //0.0625pi/1024
   sin[321]  =  14'b00001100100001;     //0.062695pi/1024
   cos[321]  =  14'b00111110110000;     //0.062695pi/1024
   sin[322]  =  14'b00001100100100;     //0.062891pi/1024
   cos[322]  =  14'b00111110110000;     //0.062891pi/1024
   sin[323]  =  14'b00001100100110;     //0.063086pi/1024
   cos[323]  =  14'b00111110101111;     //0.063086pi/1024
   sin[324]  =  14'b00001100101000;     //0.063281pi/1024
   cos[324]  =  14'b00111110101111;     //0.063281pi/1024
   sin[325]  =  14'b00001100101011;     //0.063477pi/1024
   cos[325]  =  14'b00111110101110;     //0.063477pi/1024
   sin[326]  =  14'b00001100101101;     //0.063672pi/1024
   cos[326]  =  14'b00111110101110;     //0.063672pi/1024
   sin[327]  =  14'b00001100110000;     //0.063867pi/1024
   cos[327]  =  14'b00111110101101;     //0.063867pi/1024
   sin[328]  =  14'b00001100110010;     //0.064063pi/1024
   cos[328]  =  14'b00111110101101;     //0.064063pi/1024
   sin[329]  =  14'b00001100110101;     //0.064258pi/1024
   cos[329]  =  14'b00111110101100;     //0.064258pi/1024
   sin[330]  =  14'b00001100110111;     //0.064453pi/1024
   cos[330]  =  14'b00111110101100;     //0.064453pi/1024
   sin[331]  =  14'b00001100111010;     //0.064648pi/1024
   cos[331]  =  14'b00111110101011;     //0.064648pi/1024
   sin[332]  =  14'b00001100111100;     //0.064844pi/1024
   cos[332]  =  14'b00111110101011;     //0.064844pi/1024
   sin[333]  =  14'b00001100111111;     //0.065039pi/1024
   cos[333]  =  14'b00111110101010;     //0.065039pi/1024
   sin[334]  =  14'b00001101000001;     //0.065234pi/1024
   cos[334]  =  14'b00111110101010;     //0.065234pi/1024
   sin[335]  =  14'b00001101000100;     //0.06543pi/1024
   cos[335]  =  14'b00111110101001;     //0.06543pi/1024
   sin[336]  =  14'b00001101000110;     //0.065625pi/1024
   cos[336]  =  14'b00111110101001;     //0.065625pi/1024
   sin[337]  =  14'b00001101001000;     //0.06582pi/1024
   cos[337]  =  14'b00111110101000;     //0.06582pi/1024
   sin[338]  =  14'b00001101001011;     //0.066016pi/1024
   cos[338]  =  14'b00111110101000;     //0.066016pi/1024
   sin[339]  =  14'b00001101001101;     //0.066211pi/1024
   cos[339]  =  14'b00111110100111;     //0.066211pi/1024
   sin[340]  =  14'b00001101010000;     //0.066406pi/1024
   cos[340]  =  14'b00111110100111;     //0.066406pi/1024
   sin[341]  =  14'b00001101010010;     //0.066602pi/1024
   cos[341]  =  14'b00111110100110;     //0.066602pi/1024
   sin[342]  =  14'b00001101010101;     //0.066797pi/1024
   cos[342]  =  14'b00111110100110;     //0.066797pi/1024
   sin[343]  =  14'b00001101010111;     //0.066992pi/1024
   cos[343]  =  14'b00111110100101;     //0.066992pi/1024
   sin[344]  =  14'b00001101011010;     //0.067187pi/1024
   cos[344]  =  14'b00111110100101;     //0.067187pi/1024
   sin[345]  =  14'b00001101011100;     //0.067383pi/1024
   cos[345]  =  14'b00111110100100;     //0.067383pi/1024
   sin[346]  =  14'b00001101011111;     //0.067578pi/1024
   cos[346]  =  14'b00111110100100;     //0.067578pi/1024
   sin[347]  =  14'b00001101100001;     //0.067773pi/1024
   cos[347]  =  14'b00111110100011;     //0.067773pi/1024
   sin[348]  =  14'b00001101100011;     //0.067969pi/1024
   cos[348]  =  14'b00111110100010;     //0.067969pi/1024
   sin[349]  =  14'b00001101100110;     //0.068164pi/1024
   cos[349]  =  14'b00111110100010;     //0.068164pi/1024
   sin[350]  =  14'b00001101101000;     //0.068359pi/1024
   cos[350]  =  14'b00111110100001;     //0.068359pi/1024
   sin[351]  =  14'b00001101101011;     //0.068555pi/1024
   cos[351]  =  14'b00111110100001;     //0.068555pi/1024
   sin[352]  =  14'b00001101101101;     //0.06875pi/1024
   cos[352]  =  14'b00111110100000;     //0.06875pi/1024
   sin[353]  =  14'b00001101110000;     //0.068945pi/1024
   cos[353]  =  14'b00111110100000;     //0.068945pi/1024
   sin[354]  =  14'b00001101110010;     //0.069141pi/1024
   cos[354]  =  14'b00111110011111;     //0.069141pi/1024
   sin[355]  =  14'b00001101110101;     //0.069336pi/1024
   cos[355]  =  14'b00111110011111;     //0.069336pi/1024
   sin[356]  =  14'b00001101110111;     //0.069531pi/1024
   cos[356]  =  14'b00111110011110;     //0.069531pi/1024
   sin[357]  =  14'b00001101111010;     //0.069727pi/1024
   cos[357]  =  14'b00111110011110;     //0.069727pi/1024
   sin[358]  =  14'b00001101111100;     //0.069922pi/1024
   cos[358]  =  14'b00111110011101;     //0.069922pi/1024
   sin[359]  =  14'b00001101111110;     //0.070117pi/1024
   cos[359]  =  14'b00111110011101;     //0.070117pi/1024
   sin[360]  =  14'b00001110000001;     //0.070312pi/1024
   cos[360]  =  14'b00111110011100;     //0.070312pi/1024
   sin[361]  =  14'b00001110000011;     //0.070508pi/1024
   cos[361]  =  14'b00111110011011;     //0.070508pi/1024
   sin[362]  =  14'b00001110000110;     //0.070703pi/1024
   cos[362]  =  14'b00111110011011;     //0.070703pi/1024
   sin[363]  =  14'b00001110001000;     //0.070898pi/1024
   cos[363]  =  14'b00111110011010;     //0.070898pi/1024
   sin[364]  =  14'b00001110001011;     //0.071094pi/1024
   cos[364]  =  14'b00111110011010;     //0.071094pi/1024
   sin[365]  =  14'b00001110001101;     //0.071289pi/1024
   cos[365]  =  14'b00111110011001;     //0.071289pi/1024
   sin[366]  =  14'b00001110010000;     //0.071484pi/1024
   cos[366]  =  14'b00111110011001;     //0.071484pi/1024
   sin[367]  =  14'b00001110010010;     //0.07168pi/1024
   cos[367]  =  14'b00111110011000;     //0.07168pi/1024
   sin[368]  =  14'b00001110010101;     //0.071875pi/1024
   cos[368]  =  14'b00111110011000;     //0.071875pi/1024
   sin[369]  =  14'b00001110010111;     //0.07207pi/1024
   cos[369]  =  14'b00111110010111;     //0.07207pi/1024
   sin[370]  =  14'b00001110011001;     //0.072266pi/1024
   cos[370]  =  14'b00111110010110;     //0.072266pi/1024
   sin[371]  =  14'b00001110011100;     //0.072461pi/1024
   cos[371]  =  14'b00111110010110;     //0.072461pi/1024
   sin[372]  =  14'b00001110011110;     //0.072656pi/1024
   cos[372]  =  14'b00111110010101;     //0.072656pi/1024
   sin[373]  =  14'b00001110100001;     //0.072852pi/1024
   cos[373]  =  14'b00111110010101;     //0.072852pi/1024
   sin[374]  =  14'b00001110100011;     //0.073047pi/1024
   cos[374]  =  14'b00111110010100;     //0.073047pi/1024
   sin[375]  =  14'b00001110100110;     //0.073242pi/1024
   cos[375]  =  14'b00111110010100;     //0.073242pi/1024
   sin[376]  =  14'b00001110101000;     //0.073438pi/1024
   cos[376]  =  14'b00111110010011;     //0.073438pi/1024
   sin[377]  =  14'b00001110101011;     //0.073633pi/1024
   cos[377]  =  14'b00111110010010;     //0.073633pi/1024
   sin[378]  =  14'b00001110101101;     //0.073828pi/1024
   cos[378]  =  14'b00111110010010;     //0.073828pi/1024
   sin[379]  =  14'b00001110101111;     //0.074023pi/1024
   cos[379]  =  14'b00111110010001;     //0.074023pi/1024
   sin[380]  =  14'b00001110110010;     //0.074219pi/1024
   cos[380]  =  14'b00111110010001;     //0.074219pi/1024
   sin[381]  =  14'b00001110110100;     //0.074414pi/1024
   cos[381]  =  14'b00111110010000;     //0.074414pi/1024
   sin[382]  =  14'b00001110110111;     //0.074609pi/1024
   cos[382]  =  14'b00111110001111;     //0.074609pi/1024
   sin[383]  =  14'b00001110111001;     //0.074805pi/1024
   cos[383]  =  14'b00111110001111;     //0.074805pi/1024
   sin[384]  =  14'b00001110111100;     //0.075pi/1024
   cos[384]  =  14'b00111110001110;     //0.075pi/1024
   sin[385]  =  14'b00001110111110;     //0.075195pi/1024
   cos[385]  =  14'b00111110001110;     //0.075195pi/1024
   sin[386]  =  14'b00001111000001;     //0.075391pi/1024
   cos[386]  =  14'b00111110001101;     //0.075391pi/1024
   sin[387]  =  14'b00001111000011;     //0.075586pi/1024
   cos[387]  =  14'b00111110001101;     //0.075586pi/1024
   sin[388]  =  14'b00001111000101;     //0.075781pi/1024
   cos[388]  =  14'b00111110001100;     //0.075781pi/1024
   sin[389]  =  14'b00001111001000;     //0.075977pi/1024
   cos[389]  =  14'b00111110001011;     //0.075977pi/1024
   sin[390]  =  14'b00001111001010;     //0.076172pi/1024
   cos[390]  =  14'b00111110001011;     //0.076172pi/1024
   sin[391]  =  14'b00001111001101;     //0.076367pi/1024
   cos[391]  =  14'b00111110001010;     //0.076367pi/1024
   sin[392]  =  14'b00001111001111;     //0.076563pi/1024
   cos[392]  =  14'b00111110001010;     //0.076563pi/1024
   sin[393]  =  14'b00001111010010;     //0.076758pi/1024
   cos[393]  =  14'b00111110001001;     //0.076758pi/1024
   sin[394]  =  14'b00001111010100;     //0.076953pi/1024
   cos[394]  =  14'b00111110001000;     //0.076953pi/1024
   sin[395]  =  14'b00001111010111;     //0.077148pi/1024
   cos[395]  =  14'b00111110001000;     //0.077148pi/1024
   sin[396]  =  14'b00001111011001;     //0.077344pi/1024
   cos[396]  =  14'b00111110000111;     //0.077344pi/1024
   sin[397]  =  14'b00001111011011;     //0.077539pi/1024
   cos[397]  =  14'b00111110000111;     //0.077539pi/1024
   sin[398]  =  14'b00001111011110;     //0.077734pi/1024
   cos[398]  =  14'b00111110000110;     //0.077734pi/1024
   sin[399]  =  14'b00001111100000;     //0.07793pi/1024
   cos[399]  =  14'b00111110000101;     //0.07793pi/1024
   sin[400]  =  14'b00001111100011;     //0.078125pi/1024
   cos[400]  =  14'b00111110000101;     //0.078125pi/1024
   sin[401]  =  14'b00001111100101;     //0.07832pi/1024
   cos[401]  =  14'b00111110000100;     //0.07832pi/1024
   sin[402]  =  14'b00001111101000;     //0.078516pi/1024
   cos[402]  =  14'b00111110000100;     //0.078516pi/1024
   sin[403]  =  14'b00001111101010;     //0.078711pi/1024
   cos[403]  =  14'b00111110000011;     //0.078711pi/1024
   sin[404]  =  14'b00001111101100;     //0.078906pi/1024
   cos[404]  =  14'b00111110000010;     //0.078906pi/1024
   sin[405]  =  14'b00001111101111;     //0.079102pi/1024
   cos[405]  =  14'b00111110000010;     //0.079102pi/1024
   sin[406]  =  14'b00001111110001;     //0.079297pi/1024
   cos[406]  =  14'b00111110000001;     //0.079297pi/1024
   sin[407]  =  14'b00001111110100;     //0.079492pi/1024
   cos[407]  =  14'b00111110000000;     //0.079492pi/1024
   sin[408]  =  14'b00001111110110;     //0.079688pi/1024
   cos[408]  =  14'b00111110000000;     //0.079688pi/1024
   sin[409]  =  14'b00001111111001;     //0.079883pi/1024
   cos[409]  =  14'b00111101111111;     //0.079883pi/1024
   sin[410]  =  14'b00001111111011;     //0.080078pi/1024
   cos[410]  =  14'b00111101111111;     //0.080078pi/1024
   sin[411]  =  14'b00001111111110;     //0.080273pi/1024
   cos[411]  =  14'b00111101111110;     //0.080273pi/1024
   sin[412]  =  14'b00010000000000;     //0.080469pi/1024
   cos[412]  =  14'b00111101111101;     //0.080469pi/1024
   sin[413]  =  14'b00010000000010;     //0.080664pi/1024
   cos[413]  =  14'b00111101111101;     //0.080664pi/1024
   sin[414]  =  14'b00010000000101;     //0.080859pi/1024
   cos[414]  =  14'b00111101111100;     //0.080859pi/1024
   sin[415]  =  14'b00010000000111;     //0.081055pi/1024
   cos[415]  =  14'b00111101111011;     //0.081055pi/1024
   sin[416]  =  14'b00010000001010;     //0.08125pi/1024
   cos[416]  =  14'b00111101111011;     //0.08125pi/1024
   sin[417]  =  14'b00010000001100;     //0.081445pi/1024
   cos[417]  =  14'b00111101111010;     //0.081445pi/1024
   sin[418]  =  14'b00010000001111;     //0.081641pi/1024
   cos[418]  =  14'b00111101111010;     //0.081641pi/1024
   sin[419]  =  14'b00010000010001;     //0.081836pi/1024
   cos[419]  =  14'b00111101111001;     //0.081836pi/1024
   sin[420]  =  14'b00010000010011;     //0.082031pi/1024
   cos[420]  =  14'b00111101111000;     //0.082031pi/1024
   sin[421]  =  14'b00010000010110;     //0.082227pi/1024
   cos[421]  =  14'b00111101111000;     //0.082227pi/1024
   sin[422]  =  14'b00010000011000;     //0.082422pi/1024
   cos[422]  =  14'b00111101110111;     //0.082422pi/1024
   sin[423]  =  14'b00010000011011;     //0.082617pi/1024
   cos[423]  =  14'b00111101110110;     //0.082617pi/1024
   sin[424]  =  14'b00010000011101;     //0.082813pi/1024
   cos[424]  =  14'b00111101110110;     //0.082813pi/1024
   sin[425]  =  14'b00010000100000;     //0.083008pi/1024
   cos[425]  =  14'b00111101110101;     //0.083008pi/1024
   sin[426]  =  14'b00010000100010;     //0.083203pi/1024
   cos[426]  =  14'b00111101110100;     //0.083203pi/1024
   sin[427]  =  14'b00010000100100;     //0.083398pi/1024
   cos[427]  =  14'b00111101110100;     //0.083398pi/1024
   sin[428]  =  14'b00010000100111;     //0.083594pi/1024
   cos[428]  =  14'b00111101110011;     //0.083594pi/1024
   sin[429]  =  14'b00010000101001;     //0.083789pi/1024
   cos[429]  =  14'b00111101110010;     //0.083789pi/1024
   sin[430]  =  14'b00010000101100;     //0.083984pi/1024
   cos[430]  =  14'b00111101110010;     //0.083984pi/1024
   sin[431]  =  14'b00010000101110;     //0.08418pi/1024
   cos[431]  =  14'b00111101110001;     //0.08418pi/1024
   sin[432]  =  14'b00010000110001;     //0.084375pi/1024
   cos[432]  =  14'b00111101110000;     //0.084375pi/1024
   sin[433]  =  14'b00010000110011;     //0.08457pi/1024
   cos[433]  =  14'b00111101110000;     //0.08457pi/1024
   sin[434]  =  14'b00010000110101;     //0.084766pi/1024
   cos[434]  =  14'b00111101101111;     //0.084766pi/1024
   sin[435]  =  14'b00010000111000;     //0.084961pi/1024
   cos[435]  =  14'b00111101101110;     //0.084961pi/1024
   sin[436]  =  14'b00010000111010;     //0.085156pi/1024
   cos[436]  =  14'b00111101101110;     //0.085156pi/1024
   sin[437]  =  14'b00010000111101;     //0.085352pi/1024
   cos[437]  =  14'b00111101101101;     //0.085352pi/1024
   sin[438]  =  14'b00010000111111;     //0.085547pi/1024
   cos[438]  =  14'b00111101101100;     //0.085547pi/1024
   sin[439]  =  14'b00010001000010;     //0.085742pi/1024
   cos[439]  =  14'b00111101101100;     //0.085742pi/1024
   sin[440]  =  14'b00010001000100;     //0.085938pi/1024
   cos[440]  =  14'b00111101101011;     //0.085938pi/1024
   sin[441]  =  14'b00010001000110;     //0.086133pi/1024
   cos[441]  =  14'b00111101101010;     //0.086133pi/1024
   sin[442]  =  14'b00010001001001;     //0.086328pi/1024
   cos[442]  =  14'b00111101101010;     //0.086328pi/1024
   sin[443]  =  14'b00010001001011;     //0.086523pi/1024
   cos[443]  =  14'b00111101101001;     //0.086523pi/1024
   sin[444]  =  14'b00010001001110;     //0.086719pi/1024
   cos[444]  =  14'b00111101101000;     //0.086719pi/1024
   sin[445]  =  14'b00010001010000;     //0.086914pi/1024
   cos[445]  =  14'b00111101101000;     //0.086914pi/1024
   sin[446]  =  14'b00010001010010;     //0.087109pi/1024
   cos[446]  =  14'b00111101100111;     //0.087109pi/1024
   sin[447]  =  14'b00010001010101;     //0.087305pi/1024
   cos[447]  =  14'b00111101100110;     //0.087305pi/1024
   sin[448]  =  14'b00010001010111;     //0.0875pi/1024
   cos[448]  =  14'b00111101100110;     //0.0875pi/1024
   sin[449]  =  14'b00010001011010;     //0.087695pi/1024
   cos[449]  =  14'b00111101100101;     //0.087695pi/1024
   sin[450]  =  14'b00010001011100;     //0.087891pi/1024
   cos[450]  =  14'b00111101100100;     //0.087891pi/1024
   sin[451]  =  14'b00010001011111;     //0.088086pi/1024
   cos[451]  =  14'b00111101100100;     //0.088086pi/1024
   sin[452]  =  14'b00010001100001;     //0.088281pi/1024
   cos[452]  =  14'b00111101100011;     //0.088281pi/1024
   sin[453]  =  14'b00010001100011;     //0.088477pi/1024
   cos[453]  =  14'b00111101100010;     //0.088477pi/1024
   sin[454]  =  14'b00010001100110;     //0.088672pi/1024
   cos[454]  =  14'b00111101100010;     //0.088672pi/1024
   sin[455]  =  14'b00010001101000;     //0.088867pi/1024
   cos[455]  =  14'b00111101100001;     //0.088867pi/1024
   sin[456]  =  14'b00010001101011;     //0.089063pi/1024
   cos[456]  =  14'b00111101100000;     //0.089063pi/1024
   sin[457]  =  14'b00010001101101;     //0.089258pi/1024
   cos[457]  =  14'b00111101100000;     //0.089258pi/1024
   sin[458]  =  14'b00010001101111;     //0.089453pi/1024
   cos[458]  =  14'b00111101011111;     //0.089453pi/1024
   sin[459]  =  14'b00010001110010;     //0.089648pi/1024
   cos[459]  =  14'b00111101011110;     //0.089648pi/1024
   sin[460]  =  14'b00010001110100;     //0.089844pi/1024
   cos[460]  =  14'b00111101011101;     //0.089844pi/1024
   sin[461]  =  14'b00010001110111;     //0.090039pi/1024
   cos[461]  =  14'b00111101011101;     //0.090039pi/1024
   sin[462]  =  14'b00010001111001;     //0.090234pi/1024
   cos[462]  =  14'b00111101011100;     //0.090234pi/1024
   sin[463]  =  14'b00010001111100;     //0.09043pi/1024
   cos[463]  =  14'b00111101011011;     //0.09043pi/1024
   sin[464]  =  14'b00010001111110;     //0.090625pi/1024
   cos[464]  =  14'b00111101011011;     //0.090625pi/1024
   sin[465]  =  14'b00010010000000;     //0.09082pi/1024
   cos[465]  =  14'b00111101011010;     //0.09082pi/1024
   sin[466]  =  14'b00010010000011;     //0.091016pi/1024
   cos[466]  =  14'b00111101011001;     //0.091016pi/1024
   sin[467]  =  14'b00010010000101;     //0.091211pi/1024
   cos[467]  =  14'b00111101011000;     //0.091211pi/1024
   sin[468]  =  14'b00010010001000;     //0.091406pi/1024
   cos[468]  =  14'b00111101011000;     //0.091406pi/1024
   sin[469]  =  14'b00010010001010;     //0.091602pi/1024
   cos[469]  =  14'b00111101010111;     //0.091602pi/1024
   sin[470]  =  14'b00010010001100;     //0.091797pi/1024
   cos[470]  =  14'b00111101010110;     //0.091797pi/1024
   sin[471]  =  14'b00010010001111;     //0.091992pi/1024
   cos[471]  =  14'b00111101010110;     //0.091992pi/1024
   sin[472]  =  14'b00010010010001;     //0.092188pi/1024
   cos[472]  =  14'b00111101010101;     //0.092188pi/1024
   sin[473]  =  14'b00010010010100;     //0.092383pi/1024
   cos[473]  =  14'b00111101010100;     //0.092383pi/1024
   sin[474]  =  14'b00010010010110;     //0.092578pi/1024
   cos[474]  =  14'b00111101010011;     //0.092578pi/1024
   sin[475]  =  14'b00010010011000;     //0.092773pi/1024
   cos[475]  =  14'b00111101010011;     //0.092773pi/1024
   sin[476]  =  14'b00010010011011;     //0.092969pi/1024
   cos[476]  =  14'b00111101010010;     //0.092969pi/1024
   sin[477]  =  14'b00010010011101;     //0.093164pi/1024
   cos[477]  =  14'b00111101010001;     //0.093164pi/1024
   sin[478]  =  14'b00010010100000;     //0.093359pi/1024
   cos[478]  =  14'b00111101010001;     //0.093359pi/1024
   sin[479]  =  14'b00010010100010;     //0.093555pi/1024
   cos[479]  =  14'b00111101010000;     //0.093555pi/1024
   sin[480]  =  14'b00010010100101;     //0.09375pi/1024
   cos[480]  =  14'b00111101001111;     //0.09375pi/1024
   sin[481]  =  14'b00010010100111;     //0.093945pi/1024
   cos[481]  =  14'b00111101001110;     //0.093945pi/1024
   sin[482]  =  14'b00010010101001;     //0.094141pi/1024
   cos[482]  =  14'b00111101001110;     //0.094141pi/1024
   sin[483]  =  14'b00010010101100;     //0.094336pi/1024
   cos[483]  =  14'b00111101001101;     //0.094336pi/1024
   sin[484]  =  14'b00010010101110;     //0.094531pi/1024
   cos[484]  =  14'b00111101001100;     //0.094531pi/1024
   sin[485]  =  14'b00010010110001;     //0.094727pi/1024
   cos[485]  =  14'b00111101001011;     //0.094727pi/1024
   sin[486]  =  14'b00010010110011;     //0.094922pi/1024
   cos[486]  =  14'b00111101001011;     //0.094922pi/1024
   sin[487]  =  14'b00010010110101;     //0.095117pi/1024
   cos[487]  =  14'b00111101001010;     //0.095117pi/1024
   sin[488]  =  14'b00010010111000;     //0.095313pi/1024
   cos[488]  =  14'b00111101001001;     //0.095313pi/1024
   sin[489]  =  14'b00010010111010;     //0.095508pi/1024
   cos[489]  =  14'b00111101001001;     //0.095508pi/1024
   sin[490]  =  14'b00010010111101;     //0.095703pi/1024
   cos[490]  =  14'b00111101001000;     //0.095703pi/1024
   sin[491]  =  14'b00010010111111;     //0.095898pi/1024
   cos[491]  =  14'b00111101000111;     //0.095898pi/1024
   sin[492]  =  14'b00010011000001;     //0.096094pi/1024
   cos[492]  =  14'b00111101000110;     //0.096094pi/1024
   sin[493]  =  14'b00010011000100;     //0.096289pi/1024
   cos[493]  =  14'b00111101000110;     //0.096289pi/1024
   sin[494]  =  14'b00010011000110;     //0.096484pi/1024
   cos[494]  =  14'b00111101000101;     //0.096484pi/1024
   sin[495]  =  14'b00010011001001;     //0.09668pi/1024
   cos[495]  =  14'b00111101000100;     //0.09668pi/1024
   sin[496]  =  14'b00010011001011;     //0.096875pi/1024
   cos[496]  =  14'b00111101000011;     //0.096875pi/1024
   sin[497]  =  14'b00010011001101;     //0.09707pi/1024
   cos[497]  =  14'b00111101000011;     //0.09707pi/1024
   sin[498]  =  14'b00010011010000;     //0.097266pi/1024
   cos[498]  =  14'b00111101000010;     //0.097266pi/1024
   sin[499]  =  14'b00010011010010;     //0.097461pi/1024
   cos[499]  =  14'b00111101000001;     //0.097461pi/1024
   sin[500]  =  14'b00010011010101;     //0.097656pi/1024
   cos[500]  =  14'b00111101000000;     //0.097656pi/1024
   sin[501]  =  14'b00010011010111;     //0.097852pi/1024
   cos[501]  =  14'b00111100111111;     //0.097852pi/1024
   sin[502]  =  14'b00010011011001;     //0.098047pi/1024
   cos[502]  =  14'b00111100111111;     //0.098047pi/1024
   sin[503]  =  14'b00010011011100;     //0.098242pi/1024
   cos[503]  =  14'b00111100111110;     //0.098242pi/1024
   sin[504]  =  14'b00010011011110;     //0.098438pi/1024
   cos[504]  =  14'b00111100111101;     //0.098438pi/1024
   sin[505]  =  14'b00010011100000;     //0.098633pi/1024
   cos[505]  =  14'b00111100111100;     //0.098633pi/1024
   sin[506]  =  14'b00010011100011;     //0.098828pi/1024
   cos[506]  =  14'b00111100111100;     //0.098828pi/1024
   sin[507]  =  14'b00010011100101;     //0.099023pi/1024
   cos[507]  =  14'b00111100111011;     //0.099023pi/1024
   sin[508]  =  14'b00010011101000;     //0.099219pi/1024
   cos[508]  =  14'b00111100111010;     //0.099219pi/1024
   sin[509]  =  14'b00010011101010;     //0.099414pi/1024
   cos[509]  =  14'b00111100111001;     //0.099414pi/1024
   sin[510]  =  14'b00010011101100;     //0.099609pi/1024
   cos[510]  =  14'b00111100111001;     //0.099609pi/1024
   sin[511]  =  14'b00010011101111;     //0.099805pi/1024
   cos[511]  =  14'b00111100111000;     //0.099805pi/1024
   sin[512]  =  14'b00010011110001;     //0.1pi/1024
   cos[512]  =  14'b00111100110111;     //0.1pi/1024
   sin[513]  =  14'b00010011110100;     //0.1002pi/1024
   cos[513]  =  14'b00111100110110;     //0.1002pi/1024
   sin[514]  =  14'b00010011110110;     //0.10039pi/1024
   cos[514]  =  14'b00111100110101;     //0.10039pi/1024
   sin[515]  =  14'b00010011111000;     //0.10059pi/1024
   cos[515]  =  14'b00111100110101;     //0.10059pi/1024
   sin[516]  =  14'b00010011111011;     //0.10078pi/1024
   cos[516]  =  14'b00111100110100;     //0.10078pi/1024
   sin[517]  =  14'b00010011111101;     //0.10098pi/1024
   cos[517]  =  14'b00111100110011;     //0.10098pi/1024
   sin[518]  =  14'b00010100000000;     //0.10117pi/1024
   cos[518]  =  14'b00111100110010;     //0.10117pi/1024
   sin[519]  =  14'b00010100000010;     //0.10137pi/1024
   cos[519]  =  14'b00111100110010;     //0.10137pi/1024
   sin[520]  =  14'b00010100000100;     //0.10156pi/1024
   cos[520]  =  14'b00111100110001;     //0.10156pi/1024
   sin[521]  =  14'b00010100000111;     //0.10176pi/1024
   cos[521]  =  14'b00111100110000;     //0.10176pi/1024
   sin[522]  =  14'b00010100001001;     //0.10195pi/1024
   cos[522]  =  14'b00111100101111;     //0.10195pi/1024
   sin[523]  =  14'b00010100001011;     //0.10215pi/1024
   cos[523]  =  14'b00111100101110;     //0.10215pi/1024
   sin[524]  =  14'b00010100001110;     //0.10234pi/1024
   cos[524]  =  14'b00111100101110;     //0.10234pi/1024
   sin[525]  =  14'b00010100010000;     //0.10254pi/1024
   cos[525]  =  14'b00111100101101;     //0.10254pi/1024
   sin[526]  =  14'b00010100010011;     //0.10273pi/1024
   cos[526]  =  14'b00111100101100;     //0.10273pi/1024
   sin[527]  =  14'b00010100010101;     //0.10293pi/1024
   cos[527]  =  14'b00111100101011;     //0.10293pi/1024
   sin[528]  =  14'b00010100010111;     //0.10313pi/1024
   cos[528]  =  14'b00111100101010;     //0.10313pi/1024
   sin[529]  =  14'b00010100011010;     //0.10332pi/1024
   cos[529]  =  14'b00111100101010;     //0.10332pi/1024
   sin[530]  =  14'b00010100011100;     //0.10352pi/1024
   cos[530]  =  14'b00111100101001;     //0.10352pi/1024
   sin[531]  =  14'b00010100011111;     //0.10371pi/1024
   cos[531]  =  14'b00111100101000;     //0.10371pi/1024
   sin[532]  =  14'b00010100100001;     //0.10391pi/1024
   cos[532]  =  14'b00111100100111;     //0.10391pi/1024
   sin[533]  =  14'b00010100100011;     //0.1041pi/1024
   cos[533]  =  14'b00111100100110;     //0.1041pi/1024
   sin[534]  =  14'b00010100100110;     //0.1043pi/1024
   cos[534]  =  14'b00111100100110;     //0.1043pi/1024
   sin[535]  =  14'b00010100101000;     //0.10449pi/1024
   cos[535]  =  14'b00111100100101;     //0.10449pi/1024
   sin[536]  =  14'b00010100101010;     //0.10469pi/1024
   cos[536]  =  14'b00111100100100;     //0.10469pi/1024
   sin[537]  =  14'b00010100101101;     //0.10488pi/1024
   cos[537]  =  14'b00111100100011;     //0.10488pi/1024
   sin[538]  =  14'b00010100101111;     //0.10508pi/1024
   cos[538]  =  14'b00111100100010;     //0.10508pi/1024
   sin[539]  =  14'b00010100110010;     //0.10527pi/1024
   cos[539]  =  14'b00111100100010;     //0.10527pi/1024
   sin[540]  =  14'b00010100110100;     //0.10547pi/1024
   cos[540]  =  14'b00111100100001;     //0.10547pi/1024
   sin[541]  =  14'b00010100110110;     //0.10566pi/1024
   cos[541]  =  14'b00111100100000;     //0.10566pi/1024
   sin[542]  =  14'b00010100111001;     //0.10586pi/1024
   cos[542]  =  14'b00111100011111;     //0.10586pi/1024
   sin[543]  =  14'b00010100111011;     //0.10605pi/1024
   cos[543]  =  14'b00111100011110;     //0.10605pi/1024
   sin[544]  =  14'b00010100111101;     //0.10625pi/1024
   cos[544]  =  14'b00111100011101;     //0.10625pi/1024
   sin[545]  =  14'b00010101000000;     //0.10645pi/1024
   cos[545]  =  14'b00111100011101;     //0.10645pi/1024
   sin[546]  =  14'b00010101000010;     //0.10664pi/1024
   cos[546]  =  14'b00111100011100;     //0.10664pi/1024
   sin[547]  =  14'b00010101000101;     //0.10684pi/1024
   cos[547]  =  14'b00111100011011;     //0.10684pi/1024
   sin[548]  =  14'b00010101000111;     //0.10703pi/1024
   cos[548]  =  14'b00111100011010;     //0.10703pi/1024
   sin[549]  =  14'b00010101001001;     //0.10723pi/1024
   cos[549]  =  14'b00111100011001;     //0.10723pi/1024
   sin[550]  =  14'b00010101001100;     //0.10742pi/1024
   cos[550]  =  14'b00111100011000;     //0.10742pi/1024
   sin[551]  =  14'b00010101001110;     //0.10762pi/1024
   cos[551]  =  14'b00111100011000;     //0.10762pi/1024
   sin[552]  =  14'b00010101010000;     //0.10781pi/1024
   cos[552]  =  14'b00111100010111;     //0.10781pi/1024
   sin[553]  =  14'b00010101010011;     //0.10801pi/1024
   cos[553]  =  14'b00111100010110;     //0.10801pi/1024
   sin[554]  =  14'b00010101010101;     //0.1082pi/1024
   cos[554]  =  14'b00111100010101;     //0.1082pi/1024
   sin[555]  =  14'b00010101011000;     //0.1084pi/1024
   cos[555]  =  14'b00111100010100;     //0.1084pi/1024
   sin[556]  =  14'b00010101011010;     //0.10859pi/1024
   cos[556]  =  14'b00111100010011;     //0.10859pi/1024
   sin[557]  =  14'b00010101011100;     //0.10879pi/1024
   cos[557]  =  14'b00111100010011;     //0.10879pi/1024
   sin[558]  =  14'b00010101011111;     //0.10898pi/1024
   cos[558]  =  14'b00111100010010;     //0.10898pi/1024
   sin[559]  =  14'b00010101100001;     //0.10918pi/1024
   cos[559]  =  14'b00111100010001;     //0.10918pi/1024
   sin[560]  =  14'b00010101100011;     //0.10938pi/1024
   cos[560]  =  14'b00111100010000;     //0.10938pi/1024
   sin[561]  =  14'b00010101100110;     //0.10957pi/1024
   cos[561]  =  14'b00111100001111;     //0.10957pi/1024
   sin[562]  =  14'b00010101101000;     //0.10977pi/1024
   cos[562]  =  14'b00111100001110;     //0.10977pi/1024
   sin[563]  =  14'b00010101101010;     //0.10996pi/1024
   cos[563]  =  14'b00111100001110;     //0.10996pi/1024
   sin[564]  =  14'b00010101101101;     //0.11016pi/1024
   cos[564]  =  14'b00111100001101;     //0.11016pi/1024
   sin[565]  =  14'b00010101101111;     //0.11035pi/1024
   cos[565]  =  14'b00111100001100;     //0.11035pi/1024
   sin[566]  =  14'b00010101110010;     //0.11055pi/1024
   cos[566]  =  14'b00111100001011;     //0.11055pi/1024
   sin[567]  =  14'b00010101110100;     //0.11074pi/1024
   cos[567]  =  14'b00111100001010;     //0.11074pi/1024
   sin[568]  =  14'b00010101110110;     //0.11094pi/1024
   cos[568]  =  14'b00111100001001;     //0.11094pi/1024
   sin[569]  =  14'b00010101111001;     //0.11113pi/1024
   cos[569]  =  14'b00111100001000;     //0.11113pi/1024
   sin[570]  =  14'b00010101111011;     //0.11133pi/1024
   cos[570]  =  14'b00111100001000;     //0.11133pi/1024
   sin[571]  =  14'b00010101111101;     //0.11152pi/1024
   cos[571]  =  14'b00111100000111;     //0.11152pi/1024
   sin[572]  =  14'b00010110000000;     //0.11172pi/1024
   cos[572]  =  14'b00111100000110;     //0.11172pi/1024
   sin[573]  =  14'b00010110000010;     //0.11191pi/1024
   cos[573]  =  14'b00111100000101;     //0.11191pi/1024
   sin[574]  =  14'b00010110000100;     //0.11211pi/1024
   cos[574]  =  14'b00111100000100;     //0.11211pi/1024
   sin[575]  =  14'b00010110000111;     //0.1123pi/1024
   cos[575]  =  14'b00111100000011;     //0.1123pi/1024
   sin[576]  =  14'b00010110001001;     //0.1125pi/1024
   cos[576]  =  14'b00111100000010;     //0.1125pi/1024
   sin[577]  =  14'b00010110001100;     //0.1127pi/1024
   cos[577]  =  14'b00111100000001;     //0.1127pi/1024
   sin[578]  =  14'b00010110001110;     //0.11289pi/1024
   cos[578]  =  14'b00111100000001;     //0.11289pi/1024
   sin[579]  =  14'b00010110010000;     //0.11309pi/1024
   cos[579]  =  14'b00111100000000;     //0.11309pi/1024
   sin[580]  =  14'b00010110010011;     //0.11328pi/1024
   cos[580]  =  14'b00111011111111;     //0.11328pi/1024
   sin[581]  =  14'b00010110010101;     //0.11348pi/1024
   cos[581]  =  14'b00111011111110;     //0.11348pi/1024
   sin[582]  =  14'b00010110010111;     //0.11367pi/1024
   cos[582]  =  14'b00111011111101;     //0.11367pi/1024
   sin[583]  =  14'b00010110011010;     //0.11387pi/1024
   cos[583]  =  14'b00111011111100;     //0.11387pi/1024
   sin[584]  =  14'b00010110011100;     //0.11406pi/1024
   cos[584]  =  14'b00111011111011;     //0.11406pi/1024
   sin[585]  =  14'b00010110011110;     //0.11426pi/1024
   cos[585]  =  14'b00111011111010;     //0.11426pi/1024
   sin[586]  =  14'b00010110100001;     //0.11445pi/1024
   cos[586]  =  14'b00111011111010;     //0.11445pi/1024
   sin[587]  =  14'b00010110100011;     //0.11465pi/1024
   cos[587]  =  14'b00111011111001;     //0.11465pi/1024
   sin[588]  =  14'b00010110100101;     //0.11484pi/1024
   cos[588]  =  14'b00111011111000;     //0.11484pi/1024
   sin[589]  =  14'b00010110101000;     //0.11504pi/1024
   cos[589]  =  14'b00111011110111;     //0.11504pi/1024
   sin[590]  =  14'b00010110101010;     //0.11523pi/1024
   cos[590]  =  14'b00111011110110;     //0.11523pi/1024
   sin[591]  =  14'b00010110101101;     //0.11543pi/1024
   cos[591]  =  14'b00111011110101;     //0.11543pi/1024
   sin[592]  =  14'b00010110101111;     //0.11563pi/1024
   cos[592]  =  14'b00111011110100;     //0.11563pi/1024
   sin[593]  =  14'b00010110110001;     //0.11582pi/1024
   cos[593]  =  14'b00111011110011;     //0.11582pi/1024
   sin[594]  =  14'b00010110110100;     //0.11602pi/1024
   cos[594]  =  14'b00111011110010;     //0.11602pi/1024
   sin[595]  =  14'b00010110110110;     //0.11621pi/1024
   cos[595]  =  14'b00111011110010;     //0.11621pi/1024
   sin[596]  =  14'b00010110111000;     //0.11641pi/1024
   cos[596]  =  14'b00111011110001;     //0.11641pi/1024
   sin[597]  =  14'b00010110111011;     //0.1166pi/1024
   cos[597]  =  14'b00111011110000;     //0.1166pi/1024
   sin[598]  =  14'b00010110111101;     //0.1168pi/1024
   cos[598]  =  14'b00111011101111;     //0.1168pi/1024
   sin[599]  =  14'b00010110111111;     //0.11699pi/1024
   cos[599]  =  14'b00111011101110;     //0.11699pi/1024
   sin[600]  =  14'b00010111000010;     //0.11719pi/1024
   cos[600]  =  14'b00111011101101;     //0.11719pi/1024
   sin[601]  =  14'b00010111000100;     //0.11738pi/1024
   cos[601]  =  14'b00111011101100;     //0.11738pi/1024
   sin[602]  =  14'b00010111000110;     //0.11758pi/1024
   cos[602]  =  14'b00111011101011;     //0.11758pi/1024
   sin[603]  =  14'b00010111001001;     //0.11777pi/1024
   cos[603]  =  14'b00111011101010;     //0.11777pi/1024
   sin[604]  =  14'b00010111001011;     //0.11797pi/1024
   cos[604]  =  14'b00111011101001;     //0.11797pi/1024
   sin[605]  =  14'b00010111001101;     //0.11816pi/1024
   cos[605]  =  14'b00111011101000;     //0.11816pi/1024
   sin[606]  =  14'b00010111010000;     //0.11836pi/1024
   cos[606]  =  14'b00111011101000;     //0.11836pi/1024
   sin[607]  =  14'b00010111010010;     //0.11855pi/1024
   cos[607]  =  14'b00111011100111;     //0.11855pi/1024
   sin[608]  =  14'b00010111010100;     //0.11875pi/1024
   cos[608]  =  14'b00111011100110;     //0.11875pi/1024
   sin[609]  =  14'b00010111010111;     //0.11895pi/1024
   cos[609]  =  14'b00111011100101;     //0.11895pi/1024
   sin[610]  =  14'b00010111011001;     //0.11914pi/1024
   cos[610]  =  14'b00111011100100;     //0.11914pi/1024
   sin[611]  =  14'b00010111011011;     //0.11934pi/1024
   cos[611]  =  14'b00111011100011;     //0.11934pi/1024
   sin[612]  =  14'b00010111011110;     //0.11953pi/1024
   cos[612]  =  14'b00111011100010;     //0.11953pi/1024
   sin[613]  =  14'b00010111100000;     //0.11973pi/1024
   cos[613]  =  14'b00111011100001;     //0.11973pi/1024
   sin[614]  =  14'b00010111100010;     //0.11992pi/1024
   cos[614]  =  14'b00111011100000;     //0.11992pi/1024
   sin[615]  =  14'b00010111100101;     //0.12012pi/1024
   cos[615]  =  14'b00111011011111;     //0.12012pi/1024
   sin[616]  =  14'b00010111100111;     //0.12031pi/1024
   cos[616]  =  14'b00111011011110;     //0.12031pi/1024
   sin[617]  =  14'b00010111101001;     //0.12051pi/1024
   cos[617]  =  14'b00111011011101;     //0.12051pi/1024
   sin[618]  =  14'b00010111101100;     //0.1207pi/1024
   cos[618]  =  14'b00111011011101;     //0.1207pi/1024
   sin[619]  =  14'b00010111101110;     //0.1209pi/1024
   cos[619]  =  14'b00111011011100;     //0.1209pi/1024
   sin[620]  =  14'b00010111110000;     //0.12109pi/1024
   cos[620]  =  14'b00111011011011;     //0.12109pi/1024
   sin[621]  =  14'b00010111110011;     //0.12129pi/1024
   cos[621]  =  14'b00111011011010;     //0.12129pi/1024
   sin[622]  =  14'b00010111110101;     //0.12148pi/1024
   cos[622]  =  14'b00111011011001;     //0.12148pi/1024
   sin[623]  =  14'b00010111110111;     //0.12168pi/1024
   cos[623]  =  14'b00111011011000;     //0.12168pi/1024
   sin[624]  =  14'b00010111111010;     //0.12188pi/1024
   cos[624]  =  14'b00111011010111;     //0.12188pi/1024
   sin[625]  =  14'b00010111111100;     //0.12207pi/1024
   cos[625]  =  14'b00111011010110;     //0.12207pi/1024
   sin[626]  =  14'b00010111111110;     //0.12227pi/1024
   cos[626]  =  14'b00111011010101;     //0.12227pi/1024
   sin[627]  =  14'b00011000000001;     //0.12246pi/1024
   cos[627]  =  14'b00111011010100;     //0.12246pi/1024
   sin[628]  =  14'b00011000000011;     //0.12266pi/1024
   cos[628]  =  14'b00111011010011;     //0.12266pi/1024
   sin[629]  =  14'b00011000000101;     //0.12285pi/1024
   cos[629]  =  14'b00111011010010;     //0.12285pi/1024
   sin[630]  =  14'b00011000001000;     //0.12305pi/1024
   cos[630]  =  14'b00111011010001;     //0.12305pi/1024
   sin[631]  =  14'b00011000001010;     //0.12324pi/1024
   cos[631]  =  14'b00111011010000;     //0.12324pi/1024
   sin[632]  =  14'b00011000001100;     //0.12344pi/1024
   cos[632]  =  14'b00111011001111;     //0.12344pi/1024
   sin[633]  =  14'b00011000001111;     //0.12363pi/1024
   cos[633]  =  14'b00111011001110;     //0.12363pi/1024
   sin[634]  =  14'b00011000010001;     //0.12383pi/1024
   cos[634]  =  14'b00111011001101;     //0.12383pi/1024
   sin[635]  =  14'b00011000010011;     //0.12402pi/1024
   cos[635]  =  14'b00111011001101;     //0.12402pi/1024
   sin[636]  =  14'b00011000010110;     //0.12422pi/1024
   cos[636]  =  14'b00111011001100;     //0.12422pi/1024
   sin[637]  =  14'b00011000011000;     //0.12441pi/1024
   cos[637]  =  14'b00111011001011;     //0.12441pi/1024
   sin[638]  =  14'b00011000011010;     //0.12461pi/1024
   cos[638]  =  14'b00111011001010;     //0.12461pi/1024
   sin[639]  =  14'b00011000011101;     //0.1248pi/1024
   cos[639]  =  14'b00111011001001;     //0.1248pi/1024
   sin[640]  =  14'b00011000011111;     //0.125pi/1024
   cos[640]  =  14'b00111011001000;     //0.125pi/1024
   sin[641]  =  14'b00011000100001;     //0.1252pi/1024
   cos[641]  =  14'b00111011000111;     //0.1252pi/1024
   sin[642]  =  14'b00011000100100;     //0.12539pi/1024
   cos[642]  =  14'b00111011000110;     //0.12539pi/1024
   sin[643]  =  14'b00011000100110;     //0.12559pi/1024
   cos[643]  =  14'b00111011000101;     //0.12559pi/1024
   sin[644]  =  14'b00011000101000;     //0.12578pi/1024
   cos[644]  =  14'b00111011000100;     //0.12578pi/1024
   sin[645]  =  14'b00011000101011;     //0.12598pi/1024
   cos[645]  =  14'b00111011000011;     //0.12598pi/1024
   sin[646]  =  14'b00011000101101;     //0.12617pi/1024
   cos[646]  =  14'b00111011000010;     //0.12617pi/1024
   sin[647]  =  14'b00011000101111;     //0.12637pi/1024
   cos[647]  =  14'b00111011000001;     //0.12637pi/1024
   sin[648]  =  14'b00011000110010;     //0.12656pi/1024
   cos[648]  =  14'b00111011000000;     //0.12656pi/1024
   sin[649]  =  14'b00011000110100;     //0.12676pi/1024
   cos[649]  =  14'b00111010111111;     //0.12676pi/1024
   sin[650]  =  14'b00011000110110;     //0.12695pi/1024
   cos[650]  =  14'b00111010111110;     //0.12695pi/1024
   sin[651]  =  14'b00011000111000;     //0.12715pi/1024
   cos[651]  =  14'b00111010111101;     //0.12715pi/1024
   sin[652]  =  14'b00011000111011;     //0.12734pi/1024
   cos[652]  =  14'b00111010111100;     //0.12734pi/1024
   sin[653]  =  14'b00011000111101;     //0.12754pi/1024
   cos[653]  =  14'b00111010111011;     //0.12754pi/1024
   sin[654]  =  14'b00011000111111;     //0.12773pi/1024
   cos[654]  =  14'b00111010111010;     //0.12773pi/1024
   sin[655]  =  14'b00011001000010;     //0.12793pi/1024
   cos[655]  =  14'b00111010111001;     //0.12793pi/1024
   sin[656]  =  14'b00011001000100;     //0.12813pi/1024
   cos[656]  =  14'b00111010111000;     //0.12813pi/1024
   sin[657]  =  14'b00011001000110;     //0.12832pi/1024
   cos[657]  =  14'b00111010110111;     //0.12832pi/1024
   sin[658]  =  14'b00011001001001;     //0.12852pi/1024
   cos[658]  =  14'b00111010110110;     //0.12852pi/1024
   sin[659]  =  14'b00011001001011;     //0.12871pi/1024
   cos[659]  =  14'b00111010110101;     //0.12871pi/1024
   sin[660]  =  14'b00011001001101;     //0.12891pi/1024
   cos[660]  =  14'b00111010110100;     //0.12891pi/1024
   sin[661]  =  14'b00011001010000;     //0.1291pi/1024
   cos[661]  =  14'b00111010110011;     //0.1291pi/1024
   sin[662]  =  14'b00011001010010;     //0.1293pi/1024
   cos[662]  =  14'b00111010110010;     //0.1293pi/1024
   sin[663]  =  14'b00011001010100;     //0.12949pi/1024
   cos[663]  =  14'b00111010110001;     //0.12949pi/1024
   sin[664]  =  14'b00011001010111;     //0.12969pi/1024
   cos[664]  =  14'b00111010110000;     //0.12969pi/1024
   sin[665]  =  14'b00011001011001;     //0.12988pi/1024
   cos[665]  =  14'b00111010101111;     //0.12988pi/1024
   sin[666]  =  14'b00011001011011;     //0.13008pi/1024
   cos[666]  =  14'b00111010101110;     //0.13008pi/1024
   sin[667]  =  14'b00011001011101;     //0.13027pi/1024
   cos[667]  =  14'b00111010101101;     //0.13027pi/1024
   sin[668]  =  14'b00011001100000;     //0.13047pi/1024
   cos[668]  =  14'b00111010101100;     //0.13047pi/1024
   sin[669]  =  14'b00011001100010;     //0.13066pi/1024
   cos[669]  =  14'b00111010101011;     //0.13066pi/1024
   sin[670]  =  14'b00011001100100;     //0.13086pi/1024
   cos[670]  =  14'b00111010101010;     //0.13086pi/1024
   sin[671]  =  14'b00011001100111;     //0.13105pi/1024
   cos[671]  =  14'b00111010101001;     //0.13105pi/1024
   sin[672]  =  14'b00011001101001;     //0.13125pi/1024
   cos[672]  =  14'b00111010101000;     //0.13125pi/1024
   sin[673]  =  14'b00011001101011;     //0.13145pi/1024
   cos[673]  =  14'b00111010100111;     //0.13145pi/1024
   sin[674]  =  14'b00011001101110;     //0.13164pi/1024
   cos[674]  =  14'b00111010100110;     //0.13164pi/1024
   sin[675]  =  14'b00011001110000;     //0.13184pi/1024
   cos[675]  =  14'b00111010100101;     //0.13184pi/1024
   sin[676]  =  14'b00011001110010;     //0.13203pi/1024
   cos[676]  =  14'b00111010100100;     //0.13203pi/1024
   sin[677]  =  14'b00011001110100;     //0.13223pi/1024
   cos[677]  =  14'b00111010100011;     //0.13223pi/1024
   sin[678]  =  14'b00011001110111;     //0.13242pi/1024
   cos[678]  =  14'b00111010100010;     //0.13242pi/1024
   sin[679]  =  14'b00011001111001;     //0.13262pi/1024
   cos[679]  =  14'b00111010100001;     //0.13262pi/1024
   sin[680]  =  14'b00011001111011;     //0.13281pi/1024
   cos[680]  =  14'b00111010100000;     //0.13281pi/1024
   sin[681]  =  14'b00011001111110;     //0.13301pi/1024
   cos[681]  =  14'b00111010011111;     //0.13301pi/1024
   sin[682]  =  14'b00011010000000;     //0.1332pi/1024
   cos[682]  =  14'b00111010011110;     //0.1332pi/1024
   sin[683]  =  14'b00011010000010;     //0.1334pi/1024
   cos[683]  =  14'b00111010011101;     //0.1334pi/1024
   sin[684]  =  14'b00011010000101;     //0.13359pi/1024
   cos[684]  =  14'b00111010011100;     //0.13359pi/1024
   sin[685]  =  14'b00011010000111;     //0.13379pi/1024
   cos[685]  =  14'b00111010011011;     //0.13379pi/1024
   sin[686]  =  14'b00011010001001;     //0.13398pi/1024
   cos[686]  =  14'b00111010011010;     //0.13398pi/1024
   sin[687]  =  14'b00011010001011;     //0.13418pi/1024
   cos[687]  =  14'b00111010011001;     //0.13418pi/1024
   sin[688]  =  14'b00011010001110;     //0.13437pi/1024
   cos[688]  =  14'b00111010011000;     //0.13437pi/1024
   sin[689]  =  14'b00011010010000;     //0.13457pi/1024
   cos[689]  =  14'b00111010010111;     //0.13457pi/1024
   sin[690]  =  14'b00011010010010;     //0.13477pi/1024
   cos[690]  =  14'b00111010010110;     //0.13477pi/1024
   sin[691]  =  14'b00011010010101;     //0.13496pi/1024
   cos[691]  =  14'b00111010010101;     //0.13496pi/1024
   sin[692]  =  14'b00011010010111;     //0.13516pi/1024
   cos[692]  =  14'b00111010010100;     //0.13516pi/1024
   sin[693]  =  14'b00011010011001;     //0.13535pi/1024
   cos[693]  =  14'b00111010010011;     //0.13535pi/1024
   sin[694]  =  14'b00011010011011;     //0.13555pi/1024
   cos[694]  =  14'b00111010010010;     //0.13555pi/1024
   sin[695]  =  14'b00011010011110;     //0.13574pi/1024
   cos[695]  =  14'b00111010010001;     //0.13574pi/1024
   sin[696]  =  14'b00011010100000;     //0.13594pi/1024
   cos[696]  =  14'b00111010010000;     //0.13594pi/1024
   sin[697]  =  14'b00011010100010;     //0.13613pi/1024
   cos[697]  =  14'b00111010001111;     //0.13613pi/1024
   sin[698]  =  14'b00011010100101;     //0.13633pi/1024
   cos[698]  =  14'b00111010001110;     //0.13633pi/1024
   sin[699]  =  14'b00011010100111;     //0.13652pi/1024
   cos[699]  =  14'b00111010001100;     //0.13652pi/1024
   sin[700]  =  14'b00011010101001;     //0.13672pi/1024
   cos[700]  =  14'b00111010001011;     //0.13672pi/1024
   sin[701]  =  14'b00011010101011;     //0.13691pi/1024
   cos[701]  =  14'b00111010001010;     //0.13691pi/1024
   sin[702]  =  14'b00011010101110;     //0.13711pi/1024
   cos[702]  =  14'b00111010001001;     //0.13711pi/1024
   sin[703]  =  14'b00011010110000;     //0.1373pi/1024
   cos[703]  =  14'b00111010001000;     //0.1373pi/1024
   sin[704]  =  14'b00011010110010;     //0.1375pi/1024
   cos[704]  =  14'b00111010000111;     //0.1375pi/1024
   sin[705]  =  14'b00011010110101;     //0.1377pi/1024
   cos[705]  =  14'b00111010000110;     //0.1377pi/1024
   sin[706]  =  14'b00011010110111;     //0.13789pi/1024
   cos[706]  =  14'b00111010000101;     //0.13789pi/1024
   sin[707]  =  14'b00011010111001;     //0.13809pi/1024
   cos[707]  =  14'b00111010000100;     //0.13809pi/1024
   sin[708]  =  14'b00011010111011;     //0.13828pi/1024
   cos[708]  =  14'b00111010000011;     //0.13828pi/1024
   sin[709]  =  14'b00011010111110;     //0.13848pi/1024
   cos[709]  =  14'b00111010000010;     //0.13848pi/1024
   sin[710]  =  14'b00011011000000;     //0.13867pi/1024
   cos[710]  =  14'b00111010000001;     //0.13867pi/1024
   sin[711]  =  14'b00011011000010;     //0.13887pi/1024
   cos[711]  =  14'b00111010000000;     //0.13887pi/1024
   sin[712]  =  14'b00011011000101;     //0.13906pi/1024
   cos[712]  =  14'b00111001111111;     //0.13906pi/1024
   sin[713]  =  14'b00011011000111;     //0.13926pi/1024
   cos[713]  =  14'b00111001111110;     //0.13926pi/1024
   sin[714]  =  14'b00011011001001;     //0.13945pi/1024
   cos[714]  =  14'b00111001111101;     //0.13945pi/1024
   sin[715]  =  14'b00011011001011;     //0.13965pi/1024
   cos[715]  =  14'b00111001111100;     //0.13965pi/1024
   sin[716]  =  14'b00011011001110;     //0.13984pi/1024
   cos[716]  =  14'b00111001111011;     //0.13984pi/1024
   sin[717]  =  14'b00011011010000;     //0.14004pi/1024
   cos[717]  =  14'b00111001111001;     //0.14004pi/1024
   sin[718]  =  14'b00011011010010;     //0.14023pi/1024
   cos[718]  =  14'b00111001111000;     //0.14023pi/1024
   sin[719]  =  14'b00011011010100;     //0.14043pi/1024
   cos[719]  =  14'b00111001110111;     //0.14043pi/1024
   sin[720]  =  14'b00011011010111;     //0.14062pi/1024
   cos[720]  =  14'b00111001110110;     //0.14062pi/1024
   sin[721]  =  14'b00011011011001;     //0.14082pi/1024
   cos[721]  =  14'b00111001110101;     //0.14082pi/1024
   sin[722]  =  14'b00011011011011;     //0.14102pi/1024
   cos[722]  =  14'b00111001110100;     //0.14102pi/1024
   sin[723]  =  14'b00011011011110;     //0.14121pi/1024
   cos[723]  =  14'b00111001110011;     //0.14121pi/1024
   sin[724]  =  14'b00011011100000;     //0.14141pi/1024
   cos[724]  =  14'b00111001110010;     //0.14141pi/1024
   sin[725]  =  14'b00011011100010;     //0.1416pi/1024
   cos[725]  =  14'b00111001110001;     //0.1416pi/1024
   sin[726]  =  14'b00011011100100;     //0.1418pi/1024
   cos[726]  =  14'b00111001110000;     //0.1418pi/1024
   sin[727]  =  14'b00011011100111;     //0.14199pi/1024
   cos[727]  =  14'b00111001101111;     //0.14199pi/1024
   sin[728]  =  14'b00011011101001;     //0.14219pi/1024
   cos[728]  =  14'b00111001101110;     //0.14219pi/1024
   sin[729]  =  14'b00011011101011;     //0.14238pi/1024
   cos[729]  =  14'b00111001101101;     //0.14238pi/1024
   sin[730]  =  14'b00011011101101;     //0.14258pi/1024
   cos[730]  =  14'b00111001101011;     //0.14258pi/1024
   sin[731]  =  14'b00011011110000;     //0.14277pi/1024
   cos[731]  =  14'b00111001101010;     //0.14277pi/1024
   sin[732]  =  14'b00011011110010;     //0.14297pi/1024
   cos[732]  =  14'b00111001101001;     //0.14297pi/1024
   sin[733]  =  14'b00011011110100;     //0.14316pi/1024
   cos[733]  =  14'b00111001101000;     //0.14316pi/1024
   sin[734]  =  14'b00011011110111;     //0.14336pi/1024
   cos[734]  =  14'b00111001100111;     //0.14336pi/1024
   sin[735]  =  14'b00011011111001;     //0.14355pi/1024
   cos[735]  =  14'b00111001100110;     //0.14355pi/1024
   sin[736]  =  14'b00011011111011;     //0.14375pi/1024
   cos[736]  =  14'b00111001100101;     //0.14375pi/1024
   sin[737]  =  14'b00011011111101;     //0.14395pi/1024
   cos[737]  =  14'b00111001100100;     //0.14395pi/1024
   sin[738]  =  14'b00011100000000;     //0.14414pi/1024
   cos[738]  =  14'b00111001100011;     //0.14414pi/1024
   sin[739]  =  14'b00011100000010;     //0.14434pi/1024
   cos[739]  =  14'b00111001100010;     //0.14434pi/1024
   sin[740]  =  14'b00011100000100;     //0.14453pi/1024
   cos[740]  =  14'b00111001100000;     //0.14453pi/1024
   sin[741]  =  14'b00011100000110;     //0.14473pi/1024
   cos[741]  =  14'b00111001011111;     //0.14473pi/1024
   sin[742]  =  14'b00011100001001;     //0.14492pi/1024
   cos[742]  =  14'b00111001011110;     //0.14492pi/1024
   sin[743]  =  14'b00011100001011;     //0.14512pi/1024
   cos[743]  =  14'b00111001011101;     //0.14512pi/1024
   sin[744]  =  14'b00011100001101;     //0.14531pi/1024
   cos[744]  =  14'b00111001011100;     //0.14531pi/1024
   sin[745]  =  14'b00011100001111;     //0.14551pi/1024
   cos[745]  =  14'b00111001011011;     //0.14551pi/1024
   sin[746]  =  14'b00011100010010;     //0.1457pi/1024
   cos[746]  =  14'b00111001011010;     //0.1457pi/1024
   sin[747]  =  14'b00011100010100;     //0.1459pi/1024
   cos[747]  =  14'b00111001011001;     //0.1459pi/1024
   sin[748]  =  14'b00011100010110;     //0.14609pi/1024
   cos[748]  =  14'b00111001011000;     //0.14609pi/1024
   sin[749]  =  14'b00011100011000;     //0.14629pi/1024
   cos[749]  =  14'b00111001010110;     //0.14629pi/1024
   sin[750]  =  14'b00011100011011;     //0.14648pi/1024
   cos[750]  =  14'b00111001010101;     //0.14648pi/1024
   sin[751]  =  14'b00011100011101;     //0.14668pi/1024
   cos[751]  =  14'b00111001010100;     //0.14668pi/1024
   sin[752]  =  14'b00011100011111;     //0.14688pi/1024
   cos[752]  =  14'b00111001010011;     //0.14688pi/1024
   sin[753]  =  14'b00011100100001;     //0.14707pi/1024
   cos[753]  =  14'b00111001010010;     //0.14707pi/1024
   sin[754]  =  14'b00011100100100;     //0.14727pi/1024
   cos[754]  =  14'b00111001010001;     //0.14727pi/1024
   sin[755]  =  14'b00011100100110;     //0.14746pi/1024
   cos[755]  =  14'b00111001010000;     //0.14746pi/1024
   sin[756]  =  14'b00011100101000;     //0.14766pi/1024
   cos[756]  =  14'b00111001001111;     //0.14766pi/1024
   sin[757]  =  14'b00011100101010;     //0.14785pi/1024
   cos[757]  =  14'b00111001001110;     //0.14785pi/1024
   sin[758]  =  14'b00011100101101;     //0.14805pi/1024
   cos[758]  =  14'b00111001001100;     //0.14805pi/1024
   sin[759]  =  14'b00011100101111;     //0.14824pi/1024
   cos[759]  =  14'b00111001001011;     //0.14824pi/1024
   sin[760]  =  14'b00011100110001;     //0.14844pi/1024
   cos[760]  =  14'b00111001001010;     //0.14844pi/1024
   sin[761]  =  14'b00011100110011;     //0.14863pi/1024
   cos[761]  =  14'b00111001001001;     //0.14863pi/1024
   sin[762]  =  14'b00011100110110;     //0.14883pi/1024
   cos[762]  =  14'b00111001001000;     //0.14883pi/1024
   sin[763]  =  14'b00011100111000;     //0.14902pi/1024
   cos[763]  =  14'b00111001000111;     //0.14902pi/1024
   sin[764]  =  14'b00011100111010;     //0.14922pi/1024
   cos[764]  =  14'b00111001000110;     //0.14922pi/1024
   sin[765]  =  14'b00011100111100;     //0.14941pi/1024
   cos[765]  =  14'b00111001000100;     //0.14941pi/1024
   sin[766]  =  14'b00011100111111;     //0.14961pi/1024
   cos[766]  =  14'b00111001000011;     //0.14961pi/1024
   sin[767]  =  14'b00011101000001;     //0.1498pi/1024
   cos[767]  =  14'b00111001000010;     //0.1498pi/1024
   sin[768]  =  14'b00011101000011;     //0.15pi/1024
   cos[768]  =  14'b00111001000001;     //0.15pi/1024
   sin[769]  =  14'b00011101000101;     //0.1502pi/1024
   cos[769]  =  14'b00111001000000;     //0.1502pi/1024
   sin[770]  =  14'b00011101001000;     //0.15039pi/1024
   cos[770]  =  14'b00111000111111;     //0.15039pi/1024
   sin[771]  =  14'b00011101001010;     //0.15059pi/1024
   cos[771]  =  14'b00111000111110;     //0.15059pi/1024
   sin[772]  =  14'b00011101001100;     //0.15078pi/1024
   cos[772]  =  14'b00111000111100;     //0.15078pi/1024
   sin[773]  =  14'b00011101001110;     //0.15098pi/1024
   cos[773]  =  14'b00111000111011;     //0.15098pi/1024
   sin[774]  =  14'b00011101010000;     //0.15117pi/1024
   cos[774]  =  14'b00111000111010;     //0.15117pi/1024
   sin[775]  =  14'b00011101010011;     //0.15137pi/1024
   cos[775]  =  14'b00111000111001;     //0.15137pi/1024
   sin[776]  =  14'b00011101010101;     //0.15156pi/1024
   cos[776]  =  14'b00111000111000;     //0.15156pi/1024
   sin[777]  =  14'b00011101010111;     //0.15176pi/1024
   cos[777]  =  14'b00111000110111;     //0.15176pi/1024
   sin[778]  =  14'b00011101011001;     //0.15195pi/1024
   cos[778]  =  14'b00111000110110;     //0.15195pi/1024
   sin[779]  =  14'b00011101011100;     //0.15215pi/1024
   cos[779]  =  14'b00111000110100;     //0.15215pi/1024
   sin[780]  =  14'b00011101011110;     //0.15234pi/1024
   cos[780]  =  14'b00111000110011;     //0.15234pi/1024
   sin[781]  =  14'b00011101100000;     //0.15254pi/1024
   cos[781]  =  14'b00111000110010;     //0.15254pi/1024
   sin[782]  =  14'b00011101100010;     //0.15273pi/1024
   cos[782]  =  14'b00111000110001;     //0.15273pi/1024
   sin[783]  =  14'b00011101100101;     //0.15293pi/1024
   cos[783]  =  14'b00111000110000;     //0.15293pi/1024
   sin[784]  =  14'b00011101100111;     //0.15313pi/1024
   cos[784]  =  14'b00111000101111;     //0.15313pi/1024
   sin[785]  =  14'b00011101101001;     //0.15332pi/1024
   cos[785]  =  14'b00111000101101;     //0.15332pi/1024
   sin[786]  =  14'b00011101101011;     //0.15352pi/1024
   cos[786]  =  14'b00111000101100;     //0.15352pi/1024
   sin[787]  =  14'b00011101101101;     //0.15371pi/1024
   cos[787]  =  14'b00111000101011;     //0.15371pi/1024
   sin[788]  =  14'b00011101110000;     //0.15391pi/1024
   cos[788]  =  14'b00111000101010;     //0.15391pi/1024
   sin[789]  =  14'b00011101110010;     //0.1541pi/1024
   cos[789]  =  14'b00111000101001;     //0.1541pi/1024
   sin[790]  =  14'b00011101110100;     //0.1543pi/1024
   cos[790]  =  14'b00111000101000;     //0.1543pi/1024
   sin[791]  =  14'b00011101110110;     //0.15449pi/1024
   cos[791]  =  14'b00111000100110;     //0.15449pi/1024
   sin[792]  =  14'b00011101111001;     //0.15469pi/1024
   cos[792]  =  14'b00111000100101;     //0.15469pi/1024
   sin[793]  =  14'b00011101111011;     //0.15488pi/1024
   cos[793]  =  14'b00111000100100;     //0.15488pi/1024
   sin[794]  =  14'b00011101111101;     //0.15508pi/1024
   cos[794]  =  14'b00111000100011;     //0.15508pi/1024
   sin[795]  =  14'b00011101111111;     //0.15527pi/1024
   cos[795]  =  14'b00111000100010;     //0.15527pi/1024
   sin[796]  =  14'b00011110000001;     //0.15547pi/1024
   cos[796]  =  14'b00111000100001;     //0.15547pi/1024
   sin[797]  =  14'b00011110000100;     //0.15566pi/1024
   cos[797]  =  14'b00111000011111;     //0.15566pi/1024
   sin[798]  =  14'b00011110000110;     //0.15586pi/1024
   cos[798]  =  14'b00111000011110;     //0.15586pi/1024
   sin[799]  =  14'b00011110001000;     //0.15605pi/1024
   cos[799]  =  14'b00111000011101;     //0.15605pi/1024
   sin[800]  =  14'b00011110001010;     //0.15625pi/1024
   cos[800]  =  14'b00111000011100;     //0.15625pi/1024
   sin[801]  =  14'b00011110001101;     //0.15645pi/1024
   cos[801]  =  14'b00111000011011;     //0.15645pi/1024
   sin[802]  =  14'b00011110001111;     //0.15664pi/1024
   cos[802]  =  14'b00111000011001;     //0.15664pi/1024
   sin[803]  =  14'b00011110010001;     //0.15684pi/1024
   cos[803]  =  14'b00111000011000;     //0.15684pi/1024
   sin[804]  =  14'b00011110010011;     //0.15703pi/1024
   cos[804]  =  14'b00111000010111;     //0.15703pi/1024
   sin[805]  =  14'b00011110010101;     //0.15723pi/1024
   cos[805]  =  14'b00111000010110;     //0.15723pi/1024
   sin[806]  =  14'b00011110011000;     //0.15742pi/1024
   cos[806]  =  14'b00111000010101;     //0.15742pi/1024
   sin[807]  =  14'b00011110011010;     //0.15762pi/1024
   cos[807]  =  14'b00111000010100;     //0.15762pi/1024
   sin[808]  =  14'b00011110011100;     //0.15781pi/1024
   cos[808]  =  14'b00111000010010;     //0.15781pi/1024
   sin[809]  =  14'b00011110011110;     //0.15801pi/1024
   cos[809]  =  14'b00111000010001;     //0.15801pi/1024
   sin[810]  =  14'b00011110100000;     //0.1582pi/1024
   cos[810]  =  14'b00111000010000;     //0.1582pi/1024
   sin[811]  =  14'b00011110100011;     //0.1584pi/1024
   cos[811]  =  14'b00111000001111;     //0.1584pi/1024
   sin[812]  =  14'b00011110100101;     //0.15859pi/1024
   cos[812]  =  14'b00111000001110;     //0.15859pi/1024
   sin[813]  =  14'b00011110100111;     //0.15879pi/1024
   cos[813]  =  14'b00111000001100;     //0.15879pi/1024
   sin[814]  =  14'b00011110101001;     //0.15898pi/1024
   cos[814]  =  14'b00111000001011;     //0.15898pi/1024
   sin[815]  =  14'b00011110101100;     //0.15918pi/1024
   cos[815]  =  14'b00111000001010;     //0.15918pi/1024
   sin[816]  =  14'b00011110101110;     //0.15938pi/1024
   cos[816]  =  14'b00111000001001;     //0.15938pi/1024
   sin[817]  =  14'b00011110110000;     //0.15957pi/1024
   cos[817]  =  14'b00111000001000;     //0.15957pi/1024
   sin[818]  =  14'b00011110110010;     //0.15977pi/1024
   cos[818]  =  14'b00111000000110;     //0.15977pi/1024
   sin[819]  =  14'b00011110110100;     //0.15996pi/1024
   cos[819]  =  14'b00111000000101;     //0.15996pi/1024
   sin[820]  =  14'b00011110110111;     //0.16016pi/1024
   cos[820]  =  14'b00111000000100;     //0.16016pi/1024
   sin[821]  =  14'b00011110111001;     //0.16035pi/1024
   cos[821]  =  14'b00111000000011;     //0.16035pi/1024
   sin[822]  =  14'b00011110111011;     //0.16055pi/1024
   cos[822]  =  14'b00111000000001;     //0.16055pi/1024
   sin[823]  =  14'b00011110111101;     //0.16074pi/1024
   cos[823]  =  14'b00111000000000;     //0.16074pi/1024
   sin[824]  =  14'b00011110111111;     //0.16094pi/1024
   cos[824]  =  14'b00110111111111;     //0.16094pi/1024
   sin[825]  =  14'b00011111000010;     //0.16113pi/1024
   cos[825]  =  14'b00110111111110;     //0.16113pi/1024
   sin[826]  =  14'b00011111000100;     //0.16133pi/1024
   cos[826]  =  14'b00110111111101;     //0.16133pi/1024
   sin[827]  =  14'b00011111000110;     //0.16152pi/1024
   cos[827]  =  14'b00110111111011;     //0.16152pi/1024
   sin[828]  =  14'b00011111001000;     //0.16172pi/1024
   cos[828]  =  14'b00110111111010;     //0.16172pi/1024
   sin[829]  =  14'b00011111001010;     //0.16191pi/1024
   cos[829]  =  14'b00110111111001;     //0.16191pi/1024
   sin[830]  =  14'b00011111001101;     //0.16211pi/1024
   cos[830]  =  14'b00110111111000;     //0.16211pi/1024
   sin[831]  =  14'b00011111001111;     //0.1623pi/1024
   cos[831]  =  14'b00110111110110;     //0.1623pi/1024
   sin[832]  =  14'b00011111010001;     //0.1625pi/1024
   cos[832]  =  14'b00110111110101;     //0.1625pi/1024
   sin[833]  =  14'b00011111010011;     //0.1627pi/1024
   cos[833]  =  14'b00110111110100;     //0.1627pi/1024
   sin[834]  =  14'b00011111010101;     //0.16289pi/1024
   cos[834]  =  14'b00110111110011;     //0.16289pi/1024
   sin[835]  =  14'b00011111010111;     //0.16309pi/1024
   cos[835]  =  14'b00110111110010;     //0.16309pi/1024
   sin[836]  =  14'b00011111011010;     //0.16328pi/1024
   cos[836]  =  14'b00110111110000;     //0.16328pi/1024
   sin[837]  =  14'b00011111011100;     //0.16348pi/1024
   cos[837]  =  14'b00110111101111;     //0.16348pi/1024
   sin[838]  =  14'b00011111011110;     //0.16367pi/1024
   cos[838]  =  14'b00110111101110;     //0.16367pi/1024
   sin[839]  =  14'b00011111100000;     //0.16387pi/1024
   cos[839]  =  14'b00110111101101;     //0.16387pi/1024
   sin[840]  =  14'b00011111100010;     //0.16406pi/1024
   cos[840]  =  14'b00110111101011;     //0.16406pi/1024
   sin[841]  =  14'b00011111100101;     //0.16426pi/1024
   cos[841]  =  14'b00110111101010;     //0.16426pi/1024
   sin[842]  =  14'b00011111100111;     //0.16445pi/1024
   cos[842]  =  14'b00110111101001;     //0.16445pi/1024
   sin[843]  =  14'b00011111101001;     //0.16465pi/1024
   cos[843]  =  14'b00110111101000;     //0.16465pi/1024
   sin[844]  =  14'b00011111101011;     //0.16484pi/1024
   cos[844]  =  14'b00110111100110;     //0.16484pi/1024
   sin[845]  =  14'b00011111101101;     //0.16504pi/1024
   cos[845]  =  14'b00110111100101;     //0.16504pi/1024
   sin[846]  =  14'b00011111110000;     //0.16523pi/1024
   cos[846]  =  14'b00110111100100;     //0.16523pi/1024
   sin[847]  =  14'b00011111110010;     //0.16543pi/1024
   cos[847]  =  14'b00110111100011;     //0.16543pi/1024
   sin[848]  =  14'b00011111110100;     //0.16563pi/1024
   cos[848]  =  14'b00110111100001;     //0.16563pi/1024
   sin[849]  =  14'b00011111110110;     //0.16582pi/1024
   cos[849]  =  14'b00110111100000;     //0.16582pi/1024
   sin[850]  =  14'b00011111111000;     //0.16602pi/1024
   cos[850]  =  14'b00110111011111;     //0.16602pi/1024
   sin[851]  =  14'b00011111111010;     //0.16621pi/1024
   cos[851]  =  14'b00110111011110;     //0.16621pi/1024
   sin[852]  =  14'b00011111111101;     //0.16641pi/1024
   cos[852]  =  14'b00110111011100;     //0.16641pi/1024
   sin[853]  =  14'b00011111111111;     //0.1666pi/1024
   cos[853]  =  14'b00110111011011;     //0.1666pi/1024
   sin[854]  =  14'b00100000000001;     //0.1668pi/1024
   cos[854]  =  14'b00110111011010;     //0.1668pi/1024
   sin[855]  =  14'b00100000000011;     //0.16699pi/1024
   cos[855]  =  14'b00110111011001;     //0.16699pi/1024
   sin[856]  =  14'b00100000000101;     //0.16719pi/1024
   cos[856]  =  14'b00110111010111;     //0.16719pi/1024
   sin[857]  =  14'b00100000000111;     //0.16738pi/1024
   cos[857]  =  14'b00110111010110;     //0.16738pi/1024
   sin[858]  =  14'b00100000001010;     //0.16758pi/1024
   cos[858]  =  14'b00110111010101;     //0.16758pi/1024
   sin[859]  =  14'b00100000001100;     //0.16777pi/1024
   cos[859]  =  14'b00110111010100;     //0.16777pi/1024
   sin[860]  =  14'b00100000001110;     //0.16797pi/1024
   cos[860]  =  14'b00110111010010;     //0.16797pi/1024
   sin[861]  =  14'b00100000010000;     //0.16816pi/1024
   cos[861]  =  14'b00110111010001;     //0.16816pi/1024
   sin[862]  =  14'b00100000010010;     //0.16836pi/1024
   cos[862]  =  14'b00110111010000;     //0.16836pi/1024
   sin[863]  =  14'b00100000010101;     //0.16855pi/1024
   cos[863]  =  14'b00110111001111;     //0.16855pi/1024
   sin[864]  =  14'b00100000010111;     //0.16875pi/1024
   cos[864]  =  14'b00110111001101;     //0.16875pi/1024
   sin[865]  =  14'b00100000011001;     //0.16895pi/1024
   cos[865]  =  14'b00110111001100;     //0.16895pi/1024
   sin[866]  =  14'b00100000011011;     //0.16914pi/1024
   cos[866]  =  14'b00110111001011;     //0.16914pi/1024
   sin[867]  =  14'b00100000011101;     //0.16934pi/1024
   cos[867]  =  14'b00110111001001;     //0.16934pi/1024
   sin[868]  =  14'b00100000011111;     //0.16953pi/1024
   cos[868]  =  14'b00110111001000;     //0.16953pi/1024
   sin[869]  =  14'b00100000100010;     //0.16973pi/1024
   cos[869]  =  14'b00110111000111;     //0.16973pi/1024
   sin[870]  =  14'b00100000100100;     //0.16992pi/1024
   cos[870]  =  14'b00110111000110;     //0.16992pi/1024
   sin[871]  =  14'b00100000100110;     //0.17012pi/1024
   cos[871]  =  14'b00110111000100;     //0.17012pi/1024
   sin[872]  =  14'b00100000101000;     //0.17031pi/1024
   cos[872]  =  14'b00110111000011;     //0.17031pi/1024
   sin[873]  =  14'b00100000101010;     //0.17051pi/1024
   cos[873]  =  14'b00110111000010;     //0.17051pi/1024
   sin[874]  =  14'b00100000101100;     //0.1707pi/1024
   cos[874]  =  14'b00110111000000;     //0.1707pi/1024
   sin[875]  =  14'b00100000101110;     //0.1709pi/1024
   cos[875]  =  14'b00110110111111;     //0.1709pi/1024
   sin[876]  =  14'b00100000110001;     //0.17109pi/1024
   cos[876]  =  14'b00110110111110;     //0.17109pi/1024
   sin[877]  =  14'b00100000110011;     //0.17129pi/1024
   cos[877]  =  14'b00110110111101;     //0.17129pi/1024
   sin[878]  =  14'b00100000110101;     //0.17148pi/1024
   cos[878]  =  14'b00110110111011;     //0.17148pi/1024
   sin[879]  =  14'b00100000110111;     //0.17168pi/1024
   cos[879]  =  14'b00110110111010;     //0.17168pi/1024
   sin[880]  =  14'b00100000111001;     //0.17188pi/1024
   cos[880]  =  14'b00110110111001;     //0.17188pi/1024
   sin[881]  =  14'b00100000111011;     //0.17207pi/1024
   cos[881]  =  14'b00110110110111;     //0.17207pi/1024
   sin[882]  =  14'b00100000111110;     //0.17227pi/1024
   cos[882]  =  14'b00110110110110;     //0.17227pi/1024
   sin[883]  =  14'b00100001000000;     //0.17246pi/1024
   cos[883]  =  14'b00110110110101;     //0.17246pi/1024
   sin[884]  =  14'b00100001000010;     //0.17266pi/1024
   cos[884]  =  14'b00110110110100;     //0.17266pi/1024
   sin[885]  =  14'b00100001000100;     //0.17285pi/1024
   cos[885]  =  14'b00110110110010;     //0.17285pi/1024
   sin[886]  =  14'b00100001000110;     //0.17305pi/1024
   cos[886]  =  14'b00110110110001;     //0.17305pi/1024
   sin[887]  =  14'b00100001001000;     //0.17324pi/1024
   cos[887]  =  14'b00110110110000;     //0.17324pi/1024
   sin[888]  =  14'b00100001001010;     //0.17344pi/1024
   cos[888]  =  14'b00110110101110;     //0.17344pi/1024
   sin[889]  =  14'b00100001001101;     //0.17363pi/1024
   cos[889]  =  14'b00110110101101;     //0.17363pi/1024
   sin[890]  =  14'b00100001001111;     //0.17383pi/1024
   cos[890]  =  14'b00110110101100;     //0.17383pi/1024
   sin[891]  =  14'b00100001010001;     //0.17402pi/1024
   cos[891]  =  14'b00110110101010;     //0.17402pi/1024
   sin[892]  =  14'b00100001010011;     //0.17422pi/1024
   cos[892]  =  14'b00110110101001;     //0.17422pi/1024
   sin[893]  =  14'b00100001010101;     //0.17441pi/1024
   cos[893]  =  14'b00110110101000;     //0.17441pi/1024
   sin[894]  =  14'b00100001010111;     //0.17461pi/1024
   cos[894]  =  14'b00110110100111;     //0.17461pi/1024
   sin[895]  =  14'b00100001011010;     //0.1748pi/1024
   cos[895]  =  14'b00110110100101;     //0.1748pi/1024
   sin[896]  =  14'b00100001011100;     //0.175pi/1024
   cos[896]  =  14'b00110110100100;     //0.175pi/1024
   sin[897]  =  14'b00100001011110;     //0.1752pi/1024
   cos[897]  =  14'b00110110100011;     //0.1752pi/1024
   sin[898]  =  14'b00100001100000;     //0.17539pi/1024
   cos[898]  =  14'b00110110100001;     //0.17539pi/1024
   sin[899]  =  14'b00100001100010;     //0.17559pi/1024
   cos[899]  =  14'b00110110100000;     //0.17559pi/1024
   sin[900]  =  14'b00100001100100;     //0.17578pi/1024
   cos[900]  =  14'b00110110011111;     //0.17578pi/1024
   sin[901]  =  14'b00100001100110;     //0.17598pi/1024
   cos[901]  =  14'b00110110011101;     //0.17598pi/1024
   sin[902]  =  14'b00100001101000;     //0.17617pi/1024
   cos[902]  =  14'b00110110011100;     //0.17617pi/1024
   sin[903]  =  14'b00100001101011;     //0.17637pi/1024
   cos[903]  =  14'b00110110011011;     //0.17637pi/1024
   sin[904]  =  14'b00100001101101;     //0.17656pi/1024
   cos[904]  =  14'b00110110011001;     //0.17656pi/1024
   sin[905]  =  14'b00100001101111;     //0.17676pi/1024
   cos[905]  =  14'b00110110011000;     //0.17676pi/1024
   sin[906]  =  14'b00100001110001;     //0.17695pi/1024
   cos[906]  =  14'b00110110010111;     //0.17695pi/1024
   sin[907]  =  14'b00100001110011;     //0.17715pi/1024
   cos[907]  =  14'b00110110010101;     //0.17715pi/1024
   sin[908]  =  14'b00100001110101;     //0.17734pi/1024
   cos[908]  =  14'b00110110010100;     //0.17734pi/1024
   sin[909]  =  14'b00100001110111;     //0.17754pi/1024
   cos[909]  =  14'b00110110010011;     //0.17754pi/1024
   sin[910]  =  14'b00100001111010;     //0.17773pi/1024
   cos[910]  =  14'b00110110010001;     //0.17773pi/1024
   sin[911]  =  14'b00100001111100;     //0.17793pi/1024
   cos[911]  =  14'b00110110010000;     //0.17793pi/1024
   sin[912]  =  14'b00100001111110;     //0.17813pi/1024
   cos[912]  =  14'b00110110001111;     //0.17813pi/1024
   sin[913]  =  14'b00100010000000;     //0.17832pi/1024
   cos[913]  =  14'b00110110001101;     //0.17832pi/1024
   sin[914]  =  14'b00100010000010;     //0.17852pi/1024
   cos[914]  =  14'b00110110001100;     //0.17852pi/1024
   sin[915]  =  14'b00100010000100;     //0.17871pi/1024
   cos[915]  =  14'b00110110001011;     //0.17871pi/1024
   sin[916]  =  14'b00100010000110;     //0.17891pi/1024
   cos[916]  =  14'b00110110001001;     //0.17891pi/1024
   sin[917]  =  14'b00100010001000;     //0.1791pi/1024
   cos[917]  =  14'b00110110001000;     //0.1791pi/1024
   sin[918]  =  14'b00100010001011;     //0.1793pi/1024
   cos[918]  =  14'b00110110000111;     //0.1793pi/1024
   sin[919]  =  14'b00100010001101;     //0.17949pi/1024
   cos[919]  =  14'b00110110000101;     //0.17949pi/1024
   sin[920]  =  14'b00100010001111;     //0.17969pi/1024
   cos[920]  =  14'b00110110000100;     //0.17969pi/1024
   sin[921]  =  14'b00100010010001;     //0.17988pi/1024
   cos[921]  =  14'b00110110000011;     //0.17988pi/1024
   sin[922]  =  14'b00100010010011;     //0.18008pi/1024
   cos[922]  =  14'b00110110000001;     //0.18008pi/1024
   sin[923]  =  14'b00100010010101;     //0.18027pi/1024
   cos[923]  =  14'b00110110000000;     //0.18027pi/1024
   sin[924]  =  14'b00100010010111;     //0.18047pi/1024
   cos[924]  =  14'b00110101111111;     //0.18047pi/1024
   sin[925]  =  14'b00100010011001;     //0.18066pi/1024
   cos[925]  =  14'b00110101111101;     //0.18066pi/1024
   sin[926]  =  14'b00100010011100;     //0.18086pi/1024
   cos[926]  =  14'b00110101111100;     //0.18086pi/1024
   sin[927]  =  14'b00100010011110;     //0.18105pi/1024
   cos[927]  =  14'b00110101111011;     //0.18105pi/1024
   sin[928]  =  14'b00100010100000;     //0.18125pi/1024
   cos[928]  =  14'b00110101111001;     //0.18125pi/1024
   sin[929]  =  14'b00100010100010;     //0.18145pi/1024
   cos[929]  =  14'b00110101111000;     //0.18145pi/1024
   sin[930]  =  14'b00100010100100;     //0.18164pi/1024
   cos[930]  =  14'b00110101110111;     //0.18164pi/1024
   sin[931]  =  14'b00100010100110;     //0.18184pi/1024
   cos[931]  =  14'b00110101110101;     //0.18184pi/1024
   sin[932]  =  14'b00100010101000;     //0.18203pi/1024
   cos[932]  =  14'b00110101110100;     //0.18203pi/1024
   sin[933]  =  14'b00100010101010;     //0.18223pi/1024
   cos[933]  =  14'b00110101110010;     //0.18223pi/1024
   sin[934]  =  14'b00100010101100;     //0.18242pi/1024
   cos[934]  =  14'b00110101110001;     //0.18242pi/1024
   sin[935]  =  14'b00100010101111;     //0.18262pi/1024
   cos[935]  =  14'b00110101110000;     //0.18262pi/1024
   sin[936]  =  14'b00100010110001;     //0.18281pi/1024
   cos[936]  =  14'b00110101101110;     //0.18281pi/1024
   sin[937]  =  14'b00100010110011;     //0.18301pi/1024
   cos[937]  =  14'b00110101101101;     //0.18301pi/1024
   sin[938]  =  14'b00100010110101;     //0.1832pi/1024
   cos[938]  =  14'b00110101101100;     //0.1832pi/1024
   sin[939]  =  14'b00100010110111;     //0.1834pi/1024
   cos[939]  =  14'b00110101101010;     //0.1834pi/1024
   sin[940]  =  14'b00100010111001;     //0.18359pi/1024
   cos[940]  =  14'b00110101101001;     //0.18359pi/1024
   sin[941]  =  14'b00100010111011;     //0.18379pi/1024
   cos[941]  =  14'b00110101100111;     //0.18379pi/1024
   sin[942]  =  14'b00100010111101;     //0.18398pi/1024
   cos[942]  =  14'b00110101100110;     //0.18398pi/1024
   sin[943]  =  14'b00100010111111;     //0.18418pi/1024
   cos[943]  =  14'b00110101100101;     //0.18418pi/1024
   sin[944]  =  14'b00100011000010;     //0.18438pi/1024
   cos[944]  =  14'b00110101100011;     //0.18438pi/1024
   sin[945]  =  14'b00100011000100;     //0.18457pi/1024
   cos[945]  =  14'b00110101100010;     //0.18457pi/1024
   sin[946]  =  14'b00100011000110;     //0.18477pi/1024
   cos[946]  =  14'b00110101100001;     //0.18477pi/1024
   sin[947]  =  14'b00100011001000;     //0.18496pi/1024
   cos[947]  =  14'b00110101011111;     //0.18496pi/1024
   sin[948]  =  14'b00100011001010;     //0.18516pi/1024
   cos[948]  =  14'b00110101011110;     //0.18516pi/1024
   sin[949]  =  14'b00100011001100;     //0.18535pi/1024
   cos[949]  =  14'b00110101011100;     //0.18535pi/1024
   sin[950]  =  14'b00100011001110;     //0.18555pi/1024
   cos[950]  =  14'b00110101011011;     //0.18555pi/1024
   sin[951]  =  14'b00100011010000;     //0.18574pi/1024
   cos[951]  =  14'b00110101011010;     //0.18574pi/1024
   sin[952]  =  14'b00100011010010;     //0.18594pi/1024
   cos[952]  =  14'b00110101011000;     //0.18594pi/1024
   sin[953]  =  14'b00100011010100;     //0.18613pi/1024
   cos[953]  =  14'b00110101010111;     //0.18613pi/1024
   sin[954]  =  14'b00100011010111;     //0.18633pi/1024
   cos[954]  =  14'b00110101010110;     //0.18633pi/1024
   sin[955]  =  14'b00100011011001;     //0.18652pi/1024
   cos[955]  =  14'b00110101010100;     //0.18652pi/1024
   sin[956]  =  14'b00100011011011;     //0.18672pi/1024
   cos[956]  =  14'b00110101010011;     //0.18672pi/1024
   sin[957]  =  14'b00100011011101;     //0.18691pi/1024
   cos[957]  =  14'b00110101010001;     //0.18691pi/1024
   sin[958]  =  14'b00100011011111;     //0.18711pi/1024
   cos[958]  =  14'b00110101010000;     //0.18711pi/1024
   sin[959]  =  14'b00100011100001;     //0.1873pi/1024
   cos[959]  =  14'b00110101001111;     //0.1873pi/1024
   sin[960]  =  14'b00100011100011;     //0.1875pi/1024
   cos[960]  =  14'b00110101001101;     //0.1875pi/1024
   sin[961]  =  14'b00100011100101;     //0.1877pi/1024
   cos[961]  =  14'b00110101001100;     //0.1877pi/1024
   sin[962]  =  14'b00100011100111;     //0.18789pi/1024
   cos[962]  =  14'b00110101001010;     //0.18789pi/1024
   sin[963]  =  14'b00100011101001;     //0.18809pi/1024
   cos[963]  =  14'b00110101001001;     //0.18809pi/1024
   sin[964]  =  14'b00100011101011;     //0.18828pi/1024
   cos[964]  =  14'b00110101001000;     //0.18828pi/1024
   sin[965]  =  14'b00100011101110;     //0.18848pi/1024
   cos[965]  =  14'b00110101000110;     //0.18848pi/1024
   sin[966]  =  14'b00100011110000;     //0.18867pi/1024
   cos[966]  =  14'b00110101000101;     //0.18867pi/1024
   sin[967]  =  14'b00100011110010;     //0.18887pi/1024
   cos[967]  =  14'b00110101000011;     //0.18887pi/1024
   sin[968]  =  14'b00100011110100;     //0.18906pi/1024
   cos[968]  =  14'b00110101000010;     //0.18906pi/1024
   sin[969]  =  14'b00100011110110;     //0.18926pi/1024
   cos[969]  =  14'b00110101000001;     //0.18926pi/1024
   sin[970]  =  14'b00100011111000;     //0.18945pi/1024
   cos[970]  =  14'b00110100111111;     //0.18945pi/1024
   sin[971]  =  14'b00100011111010;     //0.18965pi/1024
   cos[971]  =  14'b00110100111110;     //0.18965pi/1024
   sin[972]  =  14'b00100011111100;     //0.18984pi/1024
   cos[972]  =  14'b00110100111100;     //0.18984pi/1024
   sin[973]  =  14'b00100011111110;     //0.19004pi/1024
   cos[973]  =  14'b00110100111011;     //0.19004pi/1024
   sin[974]  =  14'b00100100000000;     //0.19023pi/1024
   cos[974]  =  14'b00110100111010;     //0.19023pi/1024
   sin[975]  =  14'b00100100000010;     //0.19043pi/1024
   cos[975]  =  14'b00110100111000;     //0.19043pi/1024
   sin[976]  =  14'b00100100000100;     //0.19063pi/1024
   cos[976]  =  14'b00110100110111;     //0.19063pi/1024
   sin[977]  =  14'b00100100000111;     //0.19082pi/1024
   cos[977]  =  14'b00110100110101;     //0.19082pi/1024
   sin[978]  =  14'b00100100001001;     //0.19102pi/1024
   cos[978]  =  14'b00110100110100;     //0.19102pi/1024
   sin[979]  =  14'b00100100001011;     //0.19121pi/1024
   cos[979]  =  14'b00110100110010;     //0.19121pi/1024
   sin[980]  =  14'b00100100001101;     //0.19141pi/1024
   cos[980]  =  14'b00110100110001;     //0.19141pi/1024
   sin[981]  =  14'b00100100001111;     //0.1916pi/1024
   cos[981]  =  14'b00110100110000;     //0.1916pi/1024
   sin[982]  =  14'b00100100010001;     //0.1918pi/1024
   cos[982]  =  14'b00110100101110;     //0.1918pi/1024
   sin[983]  =  14'b00100100010011;     //0.19199pi/1024
   cos[983]  =  14'b00110100101101;     //0.19199pi/1024
   sin[984]  =  14'b00100100010101;     //0.19219pi/1024
   cos[984]  =  14'b00110100101011;     //0.19219pi/1024
   sin[985]  =  14'b00100100010111;     //0.19238pi/1024
   cos[985]  =  14'b00110100101010;     //0.19238pi/1024
   sin[986]  =  14'b00100100011001;     //0.19258pi/1024
   cos[986]  =  14'b00110100101000;     //0.19258pi/1024
   sin[987]  =  14'b00100100011011;     //0.19277pi/1024
   cos[987]  =  14'b00110100100111;     //0.19277pi/1024
   sin[988]  =  14'b00100100011101;     //0.19297pi/1024
   cos[988]  =  14'b00110100100110;     //0.19297pi/1024
   sin[989]  =  14'b00100100011111;     //0.19316pi/1024
   cos[989]  =  14'b00110100100100;     //0.19316pi/1024
   sin[990]  =  14'b00100100100001;     //0.19336pi/1024
   cos[990]  =  14'b00110100100011;     //0.19336pi/1024
   sin[991]  =  14'b00100100100011;     //0.19355pi/1024
   cos[991]  =  14'b00110100100001;     //0.19355pi/1024
   sin[992]  =  14'b00100100100110;     //0.19375pi/1024
   cos[992]  =  14'b00110100100000;     //0.19375pi/1024
   sin[993]  =  14'b00100100101000;     //0.19395pi/1024
   cos[993]  =  14'b00110100011110;     //0.19395pi/1024
   sin[994]  =  14'b00100100101010;     //0.19414pi/1024
   cos[994]  =  14'b00110100011101;     //0.19414pi/1024
   sin[995]  =  14'b00100100101100;     //0.19434pi/1024
   cos[995]  =  14'b00110100011100;     //0.19434pi/1024
   sin[996]  =  14'b00100100101110;     //0.19453pi/1024
   cos[996]  =  14'b00110100011010;     //0.19453pi/1024
   sin[997]  =  14'b00100100110000;     //0.19473pi/1024
   cos[997]  =  14'b00110100011001;     //0.19473pi/1024
   sin[998]  =  14'b00100100110010;     //0.19492pi/1024
   cos[998]  =  14'b00110100010111;     //0.19492pi/1024
   sin[999]  =  14'b00100100110100;     //0.19512pi/1024
   cos[999]  =  14'b00110100010110;     //0.19512pi/1024
   sin[1000]  =  14'b00100100110110;     //0.19531pi/1024
   cos[1000]  =  14'b00110100010100;     //0.19531pi/1024
   sin[1001]  =  14'b00100100111000;     //0.19551pi/1024
   cos[1001]  =  14'b00110100010011;     //0.19551pi/1024
   sin[1002]  =  14'b00100100111010;     //0.1957pi/1024
   cos[1002]  =  14'b00110100010001;     //0.1957pi/1024
   sin[1003]  =  14'b00100100111100;     //0.1959pi/1024
   cos[1003]  =  14'b00110100010000;     //0.1959pi/1024
   sin[1004]  =  14'b00100100111110;     //0.19609pi/1024
   cos[1004]  =  14'b00110100001111;     //0.19609pi/1024
   sin[1005]  =  14'b00100101000000;     //0.19629pi/1024
   cos[1005]  =  14'b00110100001101;     //0.19629pi/1024
   sin[1006]  =  14'b00100101000010;     //0.19648pi/1024
   cos[1006]  =  14'b00110100001100;     //0.19648pi/1024
   sin[1007]  =  14'b00100101000100;     //0.19668pi/1024
   cos[1007]  =  14'b00110100001010;     //0.19668pi/1024
   sin[1008]  =  14'b00100101000110;     //0.19688pi/1024
   cos[1008]  =  14'b00110100001001;     //0.19688pi/1024
   sin[1009]  =  14'b00100101001000;     //0.19707pi/1024
   cos[1009]  =  14'b00110100000111;     //0.19707pi/1024
   sin[1010]  =  14'b00100101001011;     //0.19727pi/1024
   cos[1010]  =  14'b00110100000110;     //0.19727pi/1024
   sin[1011]  =  14'b00100101001101;     //0.19746pi/1024
   cos[1011]  =  14'b00110100000100;     //0.19746pi/1024
   sin[1012]  =  14'b00100101001111;     //0.19766pi/1024
   cos[1012]  =  14'b00110100000011;     //0.19766pi/1024
   sin[1013]  =  14'b00100101010001;     //0.19785pi/1024
   cos[1013]  =  14'b00110100000001;     //0.19785pi/1024
   sin[1014]  =  14'b00100101010011;     //0.19805pi/1024
   cos[1014]  =  14'b00110100000000;     //0.19805pi/1024
   sin[1015]  =  14'b00100101010101;     //0.19824pi/1024
   cos[1015]  =  14'b00110011111110;     //0.19824pi/1024
   sin[1016]  =  14'b00100101010111;     //0.19844pi/1024
   cos[1016]  =  14'b00110011111101;     //0.19844pi/1024
   sin[1017]  =  14'b00100101011001;     //0.19863pi/1024
   cos[1017]  =  14'b00110011111100;     //0.19863pi/1024
   sin[1018]  =  14'b00100101011011;     //0.19883pi/1024
   cos[1018]  =  14'b00110011111010;     //0.19883pi/1024
   sin[1019]  =  14'b00100101011101;     //0.19902pi/1024
   cos[1019]  =  14'b00110011111001;     //0.19902pi/1024
   sin[1020]  =  14'b00100101011111;     //0.19922pi/1024
   cos[1020]  =  14'b00110011110111;     //0.19922pi/1024
   sin[1021]  =  14'b00100101100001;     //0.19941pi/1024
   cos[1021]  =  14'b00110011110110;     //0.19941pi/1024
   sin[1022]  =  14'b00100101100011;     //0.19961pi/1024
   cos[1022]  =  14'b00110011110100;     //0.19961pi/1024
   sin[1023]  =  14'b00100101100101;     //0.1998pi/1024
   cos[1023]  =  14'b00110011110011;     //0.1998pi/1024

end

endmodule