module  M_TWIDLE_8_bit #(parameter SIZE =10) (
    input            en_modify, 
    input   [10:0]   rd_ptr_angle,

    output  signed [7:0]   cos_data,
    output  signed [7:0]   sin_data
 );


wire signed [7:0]  cos  [511:0];
wire signed [7:0]  sin  [511:0];

wire signed [7:0]  cos2  [511:0];
wire signed [7:0]  sin2  [511:0];

assign cos_data =   en_modify? cos2 [rd_ptr_angle] : cos [rd_ptr_angle];
assign sin_data =   en_modify? sin2 [rd_ptr_angle] : sin [rd_ptr_angle];

  assign sin[0]  =  8'b00000000;     //0pi/512
  assign cos[0]  =  8'b01000000;     //0pi/512
  assign sin[1]  =  8'b00000000;     //1pi/512
  assign cos[1]  =  8'b00111111;     //1pi/512
  assign sin[2]  =  8'b11111111;     //2pi/512
  assign cos[2]  =  8'b00111111;     //2pi/512
  assign sin[3]  =  8'b11111111;     //3pi/512
  assign cos[3]  =  8'b00111111;     //3pi/512
  assign sin[4]  =  8'b11111110;     //4pi/512
  assign cos[4]  =  8'b00111111;     //4pi/512
  assign sin[5]  =  8'b11111110;     //5pi/512
  assign cos[5]  =  8'b00111111;     //5pi/512
  assign sin[6]  =  8'b11111110;     //6pi/512
  assign cos[6]  =  8'b00111111;     //6pi/512
  assign sin[7]  =  8'b11111101;     //7pi/512
  assign cos[7]  =  8'b00111111;     //7pi/512
  assign sin[8]  =  8'b11111101;     //8pi/512
  assign cos[8]  =  8'b00111111;     //8pi/512
  assign sin[9]  =  8'b11111100;     //9pi/512
  assign cos[9]  =  8'b00111111;     //9pi/512
  assign sin[10]  =  8'b11111100;     //10pi/512
  assign cos[10]  =  8'b00111111;     //10pi/512
  assign sin[11]  =  8'b11111100;     //11pi/512
  assign cos[11]  =  8'b00111111;     //11pi/512
  assign sin[12]  =  8'b11111011;     //12pi/512
  assign cos[12]  =  8'b00111111;     //12pi/512
  assign sin[13]  =  8'b11111011;     //13pi/512
  assign cos[13]  =  8'b00111111;     //13pi/512
  assign sin[14]  =  8'b11111011;     //14pi/512
  assign cos[14]  =  8'b00111111;     //14pi/512
  assign sin[15]  =  8'b11111010;     //15pi/512
  assign cos[15]  =  8'b00111111;     //15pi/512
  assign sin[16]  =  8'b11111010;     //16pi/512
  assign cos[16]  =  8'b00111111;     //16pi/512
  assign sin[17]  =  8'b11111001;     //17pi/512
  assign cos[17]  =  8'b00111111;     //17pi/512
  assign sin[18]  =  8'b11111001;     //18pi/512
  assign cos[18]  =  8'b00111111;     //18pi/512
  assign sin[19]  =  8'b11111001;     //19pi/512
  assign cos[19]  =  8'b00111111;     //19pi/512
  assign sin[20]  =  8'b11111000;     //20pi/512
  assign cos[20]  =  8'b00111111;     //20pi/512
  assign sin[21]  =  8'b11111000;     //21pi/512
  assign cos[21]  =  8'b00111111;     //21pi/512
  assign sin[22]  =  8'b11110111;     //22pi/512
  assign cos[22]  =  8'b00111111;     //22pi/512
  assign sin[23]  =  8'b11110111;     //23pi/512
  assign cos[23]  =  8'b00111111;     //23pi/512
  assign sin[24]  =  8'b11110111;     //24pi/512
  assign cos[24]  =  8'b00111111;     //24pi/512
  assign sin[25]  =  8'b11110110;     //25pi/512
  assign cos[25]  =  8'b00111111;     //25pi/512
  assign sin[26]  =  8'b11110110;     //26pi/512
  assign cos[26]  =  8'b00111111;     //26pi/512
  assign sin[27]  =  8'b11110101;     //27pi/512
  assign cos[27]  =  8'b00111111;     //27pi/512
  assign sin[28]  =  8'b11110101;     //28pi/512
  assign cos[28]  =  8'b00111111;     //28pi/512
  assign sin[29]  =  8'b11110101;     //29pi/512
  assign cos[29]  =  8'b00111110;     //29pi/512
  assign sin[30]  =  8'b11110100;     //30pi/512
  assign cos[30]  =  8'b00111110;     //30pi/512
  assign sin[31]  =  8'b11110100;     //31pi/512
  assign cos[31]  =  8'b00111110;     //31pi/512
  assign sin[32]  =  8'b11110100;     //32pi/512
  assign cos[32]  =  8'b00111110;     //32pi/512
  assign sin[33]  =  8'b11110011;     //33pi/512
  assign cos[33]  =  8'b00111110;     //33pi/512
  assign sin[34]  =  8'b11110011;     //34pi/512
  assign cos[34]  =  8'b00111110;     //34pi/512
  assign sin[35]  =  8'b11110010;     //35pi/512
  assign cos[35]  =  8'b00111110;     //35pi/512
  assign sin[36]  =  8'b11110010;     //36pi/512
  assign cos[36]  =  8'b00111110;     //36pi/512
  assign sin[37]  =  8'b11110010;     //37pi/512
  assign cos[37]  =  8'b00111110;     //37pi/512
  assign sin[38]  =  8'b11110001;     //38pi/512
  assign cos[38]  =  8'b00111110;     //38pi/512
  assign sin[39]  =  8'b11110001;     //39pi/512
  assign cos[39]  =  8'b00111110;     //39pi/512
  assign sin[40]  =  8'b11110000;     //40pi/512
  assign cos[40]  =  8'b00111110;     //40pi/512
  assign sin[41]  =  8'b11110000;     //41pi/512
  assign cos[41]  =  8'b00111101;     //41pi/512
  assign sin[42]  =  8'b11110000;     //42pi/512
  assign cos[42]  =  8'b00111101;     //42pi/512
  assign sin[43]  =  8'b11101111;     //43pi/512
  assign cos[43]  =  8'b00111101;     //43pi/512
  assign sin[44]  =  8'b11101111;     //44pi/512
  assign cos[44]  =  8'b00111101;     //44pi/512
  assign sin[45]  =  8'b11101111;     //45pi/512
  assign cos[45]  =  8'b00111101;     //45pi/512
  assign sin[46]  =  8'b11101110;     //46pi/512
  assign cos[46]  =  8'b00111101;     //46pi/512
  assign sin[47]  =  8'b11101110;     //47pi/512
  assign cos[47]  =  8'b00111101;     //47pi/512
  assign sin[48]  =  8'b11101101;     //48pi/512
  assign cos[48]  =  8'b00111101;     //48pi/512
  assign sin[49]  =  8'b11101101;     //49pi/512
  assign cos[49]  =  8'b00111101;     //49pi/512
  assign sin[50]  =  8'b11101101;     //50pi/512
  assign cos[50]  =  8'b00111101;     //50pi/512
  assign sin[51]  =  8'b11101100;     //51pi/512
  assign cos[51]  =  8'b00111100;     //51pi/512
  assign sin[52]  =  8'b11101100;     //52pi/512
  assign cos[52]  =  8'b00111100;     //52pi/512
  assign sin[53]  =  8'b11101100;     //53pi/512
  assign cos[53]  =  8'b00111100;     //53pi/512
  assign sin[54]  =  8'b11101011;     //54pi/512
  assign cos[54]  =  8'b00111100;     //54pi/512
  assign sin[55]  =  8'b11101011;     //55pi/512
  assign cos[55]  =  8'b00111100;     //55pi/512
  assign sin[56]  =  8'b11101010;     //56pi/512
  assign cos[56]  =  8'b00111100;     //56pi/512
  assign sin[57]  =  8'b11101010;     //57pi/512
  assign cos[57]  =  8'b00111100;     //57pi/512
  assign sin[58]  =  8'b11101010;     //58pi/512
  assign cos[58]  =  8'b00111011;     //58pi/512
  assign sin[59]  =  8'b11101001;     //59pi/512
  assign cos[59]  =  8'b00111011;     //59pi/512
  assign sin[60]  =  8'b11101001;     //60pi/512
  assign cos[60]  =  8'b00111011;     //60pi/512
  assign sin[61]  =  8'b11101001;     //61pi/512
  assign cos[61]  =  8'b00111011;     //61pi/512
  assign sin[62]  =  8'b11101000;     //62pi/512
  assign cos[62]  =  8'b00111011;     //62pi/512
  assign sin[63]  =  8'b11101000;     //63pi/512
  assign cos[63]  =  8'b00111011;     //63pi/512
  assign sin[64]  =  8'b11101000;     //64pi/512
  assign cos[64]  =  8'b00111011;     //64pi/512
  assign sin[65]  =  8'b11100111;     //65pi/512
  assign cos[65]  =  8'b00111010;     //65pi/512
  assign sin[66]  =  8'b11100111;     //66pi/512
  assign cos[66]  =  8'b00111010;     //66pi/512
  assign sin[67]  =  8'b11100110;     //67pi/512
  assign cos[67]  =  8'b00111010;     //67pi/512
  assign sin[68]  =  8'b11100110;     //68pi/512
  assign cos[68]  =  8'b00111010;     //68pi/512
  assign sin[69]  =  8'b11100110;     //69pi/512
  assign cos[69]  =  8'b00111010;     //69pi/512
  assign sin[70]  =  8'b11100101;     //70pi/512
  assign cos[70]  =  8'b00111010;     //70pi/512
  assign sin[71]  =  8'b11100101;     //71pi/512
  assign cos[71]  =  8'b00111010;     //71pi/512
  assign sin[72]  =  8'b11100101;     //72pi/512
  assign cos[72]  =  8'b00111001;     //72pi/512
  assign sin[73]  =  8'b11100100;     //73pi/512
  assign cos[73]  =  8'b00111001;     //73pi/512
  assign sin[74]  =  8'b11100100;     //74pi/512
  assign cos[74]  =  8'b00111001;     //74pi/512
  assign sin[75]  =  8'b11100100;     //75pi/512
  assign cos[75]  =  8'b00111001;     //75pi/512
  assign sin[76]  =  8'b11100011;     //76pi/512
  assign cos[76]  =  8'b00111001;     //76pi/512
  assign sin[77]  =  8'b11100011;     //77pi/512
  assign cos[77]  =  8'b00111000;     //77pi/512
  assign sin[78]  =  8'b11100011;     //78pi/512
  assign cos[78]  =  8'b00111000;     //78pi/512
  assign sin[79]  =  8'b11100010;     //79pi/512
  assign cos[79]  =  8'b00111000;     //79pi/512
  assign sin[80]  =  8'b11100010;     //80pi/512
  assign cos[80]  =  8'b00111000;     //80pi/512
  assign sin[81]  =  8'b11100001;     //81pi/512
  assign cos[81]  =  8'b00111000;     //81pi/512
  assign sin[82]  =  8'b11100001;     //82pi/512
  assign cos[82]  =  8'b00111000;     //82pi/512
  assign sin[83]  =  8'b11100001;     //83pi/512
  assign cos[83]  =  8'b00110111;     //83pi/512
  assign sin[84]  =  8'b11100000;     //84pi/512
  assign cos[84]  =  8'b00110111;     //84pi/512
  assign sin[85]  =  8'b11100000;     //85pi/512
  assign cos[85]  =  8'b00110111;     //85pi/512
  assign sin[86]  =  8'b11100000;     //86pi/512
  assign cos[86]  =  8'b00110111;     //86pi/512
  assign sin[87]  =  8'b11011111;     //87pi/512
  assign cos[87]  =  8'b00110111;     //87pi/512
  assign sin[88]  =  8'b11011111;     //88pi/512
  assign cos[88]  =  8'b00110110;     //88pi/512
  assign sin[89]  =  8'b11011111;     //89pi/512
  assign cos[89]  =  8'b00110110;     //89pi/512
  assign sin[90]  =  8'b11011110;     //90pi/512
  assign cos[90]  =  8'b00110110;     //90pi/512
  assign sin[91]  =  8'b11011110;     //91pi/512
  assign cos[91]  =  8'b00110110;     //91pi/512
  assign sin[92]  =  8'b11011110;     //92pi/512
  assign cos[92]  =  8'b00110110;     //92pi/512
  assign sin[93]  =  8'b11011101;     //93pi/512
  assign cos[93]  =  8'b00110101;     //93pi/512
  assign sin[94]  =  8'b11011101;     //94pi/512
  assign cos[94]  =  8'b00110101;     //94pi/512
  assign sin[95]  =  8'b11011101;     //95pi/512
  assign cos[95]  =  8'b00110101;     //95pi/512
  assign sin[96]  =  8'b11011100;     //96pi/512
  assign cos[96]  =  8'b00110101;     //96pi/512
  assign sin[97]  =  8'b11011100;     //97pi/512
  assign cos[97]  =  8'b00110100;     //97pi/512
  assign sin[98]  =  8'b11011100;     //98pi/512
  assign cos[98]  =  8'b00110100;     //98pi/512
  assign sin[99]  =  8'b11011011;     //99pi/512
  assign cos[99]  =  8'b00110100;     //99pi/512
  assign sin[100]  =  8'b11011011;     //100pi/512
  assign cos[100]  =  8'b00110100;     //100pi/512
  assign sin[101]  =  8'b11011011;     //101pi/512
  assign cos[101]  =  8'b00110100;     //101pi/512
  assign sin[102]  =  8'b11011011;     //102pi/512
  assign cos[102]  =  8'b00110011;     //102pi/512
  assign sin[103]  =  8'b11011010;     //103pi/512
  assign cos[103]  =  8'b00110011;     //103pi/512
  assign sin[104]  =  8'b11011010;     //104pi/512
  assign cos[104]  =  8'b00110011;     //104pi/512
  assign sin[105]  =  8'b11011010;     //105pi/512
  assign cos[105]  =  8'b00110011;     //105pi/512
  assign sin[106]  =  8'b11011001;     //106pi/512
  assign cos[106]  =  8'b00110010;     //106pi/512
  assign sin[107]  =  8'b11011001;     //107pi/512
  assign cos[107]  =  8'b00110010;     //107pi/512
  assign sin[108]  =  8'b11011001;     //108pi/512
  assign cos[108]  =  8'b00110010;     //108pi/512
  assign sin[109]  =  8'b11011000;     //109pi/512
  assign cos[109]  =  8'b00110010;     //109pi/512
  assign sin[110]  =  8'b11011000;     //110pi/512
  assign cos[110]  =  8'b00110001;     //110pi/512
  assign sin[111]  =  8'b11011000;     //111pi/512
  assign cos[111]  =  8'b00110001;     //111pi/512
  assign sin[112]  =  8'b11010111;     //112pi/512
  assign cos[112]  =  8'b00110001;     //112pi/512
  assign sin[113]  =  8'b11010111;     //113pi/512
  assign cos[113]  =  8'b00110001;     //113pi/512
  assign sin[114]  =  8'b11010111;     //114pi/512
  assign cos[114]  =  8'b00110000;     //114pi/512
  assign sin[115]  =  8'b11010110;     //115pi/512
  assign cos[115]  =  8'b00110000;     //115pi/512
  assign sin[116]  =  8'b11010110;     //116pi/512
  assign cos[116]  =  8'b00110000;     //116pi/512
  assign sin[117]  =  8'b11010110;     //117pi/512
  assign cos[117]  =  8'b00110000;     //117pi/512
  assign sin[118]  =  8'b11010110;     //118pi/512
  assign cos[118]  =  8'b00101111;     //118pi/512
  assign sin[119]  =  8'b11010101;     //119pi/512
  assign cos[119]  =  8'b00101111;     //119pi/512
  assign sin[120]  =  8'b11010101;     //120pi/512
  assign cos[120]  =  8'b00101111;     //120pi/512
  assign sin[121]  =  8'b11010101;     //121pi/512
  assign cos[121]  =  8'b00101111;     //121pi/512
  assign sin[122]  =  8'b11010100;     //122pi/512
  assign cos[122]  =  8'b00101110;     //122pi/512
  assign sin[123]  =  8'b11010100;     //123pi/512
  assign cos[123]  =  8'b00101110;     //123pi/512
  assign sin[124]  =  8'b11010100;     //124pi/512
  assign cos[124]  =  8'b00101110;     //124pi/512
  assign sin[125]  =  8'b11010100;     //125pi/512
  assign cos[125]  =  8'b00101110;     //125pi/512
  assign sin[126]  =  8'b11010011;     //126pi/512
  assign cos[126]  =  8'b00101101;     //126pi/512
  assign sin[127]  =  8'b11010011;     //127pi/512
  assign cos[127]  =  8'b00101101;     //127pi/512
  assign sin[128]  =  8'b11010011;     //128pi/512
  assign cos[128]  =  8'b00101101;     //128pi/512
  assign sin[129]  =  8'b11010010;     //129pi/512
  assign cos[129]  =  8'b00101100;     //129pi/512
  assign sin[130]  =  8'b11010010;     //130pi/512
  assign cos[130]  =  8'b00101100;     //130pi/512
  assign sin[131]  =  8'b11010010;     //131pi/512
  assign cos[131]  =  8'b00101100;     //131pi/512
  assign sin[132]  =  8'b11010010;     //132pi/512
  assign cos[132]  =  8'b00101100;     //132pi/512
  assign sin[133]  =  8'b11010001;     //133pi/512
  assign cos[133]  =  8'b00101011;     //133pi/512
  assign sin[134]  =  8'b11010001;     //134pi/512
  assign cos[134]  =  8'b00101011;     //134pi/512
  assign sin[135]  =  8'b11010001;     //135pi/512
  assign cos[135]  =  8'b00101011;     //135pi/512
  assign sin[136]  =  8'b11010001;     //136pi/512
  assign cos[136]  =  8'b00101010;     //136pi/512
  assign sin[137]  =  8'b11010000;     //137pi/512
  assign cos[137]  =  8'b00101010;     //137pi/512
  assign sin[138]  =  8'b11010000;     //138pi/512
  assign cos[138]  =  8'b00101010;     //138pi/512
  assign sin[139]  =  8'b11010000;     //139pi/512
  assign cos[139]  =  8'b00101010;     //139pi/512
  assign sin[140]  =  8'b11010000;     //140pi/512
  assign cos[140]  =  8'b00101001;     //140pi/512
  assign sin[141]  =  8'b11001111;     //141pi/512
  assign cos[141]  =  8'b00101001;     //141pi/512
  assign sin[142]  =  8'b11001111;     //142pi/512
  assign cos[142]  =  8'b00101001;     //142pi/512
  assign sin[143]  =  8'b11001111;     //143pi/512
  assign cos[143]  =  8'b00101000;     //143pi/512
  assign sin[144]  =  8'b11001111;     //144pi/512
  assign cos[144]  =  8'b00101000;     //144pi/512
  assign sin[145]  =  8'b11001110;     //145pi/512
  assign cos[145]  =  8'b00101000;     //145pi/512
  assign sin[146]  =  8'b11001110;     //146pi/512
  assign cos[146]  =  8'b00100111;     //146pi/512
  assign sin[147]  =  8'b11001110;     //147pi/512
  assign cos[147]  =  8'b00100111;     //147pi/512
  assign sin[148]  =  8'b11001110;     //148pi/512
  assign cos[148]  =  8'b00100111;     //148pi/512
  assign sin[149]  =  8'b11001101;     //149pi/512
  assign cos[149]  =  8'b00100111;     //149pi/512
  assign sin[150]  =  8'b11001101;     //150pi/512
  assign cos[150]  =  8'b00100110;     //150pi/512
  assign sin[151]  =  8'b11001101;     //151pi/512
  assign cos[151]  =  8'b00100110;     //151pi/512
  assign sin[152]  =  8'b11001101;     //152pi/512
  assign cos[152]  =  8'b00100110;     //152pi/512
  assign sin[153]  =  8'b11001100;     //153pi/512
  assign cos[153]  =  8'b00100101;     //153pi/512
  assign sin[154]  =  8'b11001100;     //154pi/512
  assign cos[154]  =  8'b00100101;     //154pi/512
  assign sin[155]  =  8'b11001100;     //155pi/512
  assign cos[155]  =  8'b00100101;     //155pi/512
  assign sin[156]  =  8'b11001100;     //156pi/512
  assign cos[156]  =  8'b00100100;     //156pi/512
  assign sin[157]  =  8'b11001011;     //157pi/512
  assign cos[157]  =  8'b00100100;     //157pi/512
  assign sin[158]  =  8'b11001011;     //158pi/512
  assign cos[158]  =  8'b00100100;     //158pi/512
  assign sin[159]  =  8'b11001011;     //159pi/512
  assign cos[159]  =  8'b00100011;     //159pi/512
  assign sin[160]  =  8'b11001011;     //160pi/512
  assign cos[160]  =  8'b00100011;     //160pi/512
  assign sin[161]  =  8'b11001011;     //161pi/512
  assign cos[161]  =  8'b00100011;     //161pi/512
  assign sin[162]  =  8'b11001010;     //162pi/512
  assign cos[162]  =  8'b00100010;     //162pi/512
  assign sin[163]  =  8'b11001010;     //163pi/512
  assign cos[163]  =  8'b00100010;     //163pi/512
  assign sin[164]  =  8'b11001010;     //164pi/512
  assign cos[164]  =  8'b00100010;     //164pi/512
  assign sin[165]  =  8'b11001010;     //165pi/512
  assign cos[165]  =  8'b00100001;     //165pi/512
  assign sin[166]  =  8'b11001010;     //166pi/512
  assign cos[166]  =  8'b00100001;     //166pi/512
  assign sin[167]  =  8'b11001001;     //167pi/512
  assign cos[167]  =  8'b00100001;     //167pi/512
  assign sin[168]  =  8'b11001001;     //168pi/512
  assign cos[168]  =  8'b00100000;     //168pi/512
  assign sin[169]  =  8'b11001001;     //169pi/512
  assign cos[169]  =  8'b00100000;     //169pi/512
  assign sin[170]  =  8'b11001001;     //170pi/512
  assign cos[170]  =  8'b00100000;     //170pi/512
  assign sin[171]  =  8'b11001001;     //171pi/512
  assign cos[171]  =  8'b00011111;     //171pi/512
  assign sin[172]  =  8'b11001000;     //172pi/512
  assign cos[172]  =  8'b00011111;     //172pi/512
  assign sin[173]  =  8'b11001000;     //173pi/512
  assign cos[173]  =  8'b00011111;     //173pi/512
  assign sin[174]  =  8'b11001000;     //174pi/512
  assign cos[174]  =  8'b00011110;     //174pi/512
  assign sin[175]  =  8'b11001000;     //175pi/512
  assign cos[175]  =  8'b00011110;     //175pi/512
  assign sin[176]  =  8'b11001000;     //176pi/512
  assign cos[176]  =  8'b00011110;     //176pi/512
  assign sin[177]  =  8'b11000111;     //177pi/512
  assign cos[177]  =  8'b00011101;     //177pi/512
  assign sin[178]  =  8'b11000111;     //178pi/512
  assign cos[178]  =  8'b00011101;     //178pi/512
  assign sin[179]  =  8'b11000111;     //179pi/512
  assign cos[179]  =  8'b00011101;     //179pi/512
  assign sin[180]  =  8'b11000111;     //180pi/512
  assign cos[180]  =  8'b00011100;     //180pi/512
  assign sin[181]  =  8'b11000111;     //181pi/512
  assign cos[181]  =  8'b00011100;     //181pi/512
  assign sin[182]  =  8'b11000110;     //182pi/512
  assign cos[182]  =  8'b00011100;     //182pi/512
  assign sin[183]  =  8'b11000110;     //183pi/512
  assign cos[183]  =  8'b00011011;     //183pi/512
  assign sin[184]  =  8'b11000110;     //184pi/512
  assign cos[184]  =  8'b00011011;     //184pi/512
  assign sin[185]  =  8'b11000110;     //185pi/512
  assign cos[185]  =  8'b00011011;     //185pi/512
  assign sin[186]  =  8'b11000110;     //186pi/512
  assign cos[186]  =  8'b00011010;     //186pi/512
  assign sin[187]  =  8'b11000110;     //187pi/512
  assign cos[187]  =  8'b00011010;     //187pi/512
  assign sin[188]  =  8'b11000101;     //188pi/512
  assign cos[188]  =  8'b00011001;     //188pi/512
  assign sin[189]  =  8'b11000101;     //189pi/512
  assign cos[189]  =  8'b00011001;     //189pi/512
  assign sin[190]  =  8'b11000101;     //190pi/512
  assign cos[190]  =  8'b00011001;     //190pi/512
  assign sin[191]  =  8'b11000101;     //191pi/512
  assign cos[191]  =  8'b00011000;     //191pi/512
  assign sin[192]  =  8'b11000101;     //192pi/512
  assign cos[192]  =  8'b00011000;     //192pi/512
  assign sin[193]  =  8'b11000101;     //193pi/512
  assign cos[193]  =  8'b00011000;     //193pi/512
  assign sin[194]  =  8'b11000101;     //194pi/512
  assign cos[194]  =  8'b00010111;     //194pi/512
  assign sin[195]  =  8'b11000100;     //195pi/512
  assign cos[195]  =  8'b00010111;     //195pi/512
  assign sin[196]  =  8'b11000100;     //196pi/512
  assign cos[196]  =  8'b00010111;     //196pi/512
  assign sin[197]  =  8'b11000100;     //197pi/512
  assign cos[197]  =  8'b00010110;     //197pi/512
  assign sin[198]  =  8'b11000100;     //198pi/512
  assign cos[198]  =  8'b00010110;     //198pi/512
  assign sin[199]  =  8'b11000100;     //199pi/512
  assign cos[199]  =  8'b00010101;     //199pi/512
  assign sin[200]  =  8'b11000100;     //200pi/512
  assign cos[200]  =  8'b00010101;     //200pi/512
  assign sin[201]  =  8'b11000100;     //201pi/512
  assign cos[201]  =  8'b00010101;     //201pi/512
  assign sin[202]  =  8'b11000011;     //202pi/512
  assign cos[202]  =  8'b00010100;     //202pi/512
  assign sin[203]  =  8'b11000011;     //203pi/512
  assign cos[203]  =  8'b00010100;     //203pi/512
  assign sin[204]  =  8'b11000011;     //204pi/512
  assign cos[204]  =  8'b00010100;     //204pi/512
  assign sin[205]  =  8'b11000011;     //205pi/512
  assign cos[205]  =  8'b00010011;     //205pi/512
  assign sin[206]  =  8'b11000011;     //206pi/512
  assign cos[206]  =  8'b00010011;     //206pi/512
  assign sin[207]  =  8'b11000011;     //207pi/512
  assign cos[207]  =  8'b00010010;     //207pi/512
  assign sin[208]  =  8'b11000011;     //208pi/512
  assign cos[208]  =  8'b00010010;     //208pi/512
  assign sin[209]  =  8'b11000011;     //209pi/512
  assign cos[209]  =  8'b00010010;     //209pi/512
  assign sin[210]  =  8'b11000011;     //210pi/512
  assign cos[210]  =  8'b00010001;     //210pi/512
  assign sin[211]  =  8'b11000010;     //211pi/512
  assign cos[211]  =  8'b00010001;     //211pi/512
  assign sin[212]  =  8'b11000010;     //212pi/512
  assign cos[212]  =  8'b00010001;     //212pi/512
  assign sin[213]  =  8'b11000010;     //213pi/512
  assign cos[213]  =  8'b00010000;     //213pi/512
  assign sin[214]  =  8'b11000010;     //214pi/512
  assign cos[214]  =  8'b00010000;     //214pi/512
  assign sin[215]  =  8'b11000010;     //215pi/512
  assign cos[215]  =  8'b00001111;     //215pi/512
  assign sin[216]  =  8'b11000010;     //216pi/512
  assign cos[216]  =  8'b00001111;     //216pi/512
  assign sin[217]  =  8'b11000010;     //217pi/512
  assign cos[217]  =  8'b00001111;     //217pi/512
  assign sin[218]  =  8'b11000010;     //218pi/512
  assign cos[218]  =  8'b00001110;     //218pi/512
  assign sin[219]  =  8'b11000010;     //219pi/512
  assign cos[219]  =  8'b00001110;     //219pi/512
  assign sin[220]  =  8'b11000010;     //220pi/512
  assign cos[220]  =  8'b00001110;     //220pi/512
  assign sin[221]  =  8'b11000001;     //221pi/512
  assign cos[221]  =  8'b00001101;     //221pi/512
  assign sin[222]  =  8'b11000001;     //222pi/512
  assign cos[222]  =  8'b00001101;     //222pi/512
  assign sin[223]  =  8'b11000001;     //223pi/512
  assign cos[223]  =  8'b00001100;     //223pi/512
  assign sin[224]  =  8'b11000001;     //224pi/512
  assign cos[224]  =  8'b00001100;     //224pi/512
  assign sin[225]  =  8'b11000001;     //225pi/512
  assign cos[225]  =  8'b00001100;     //225pi/512
  assign sin[226]  =  8'b11000001;     //226pi/512
  assign cos[226]  =  8'b00001011;     //226pi/512
  assign sin[227]  =  8'b11000001;     //227pi/512
  assign cos[227]  =  8'b00001011;     //227pi/512
  assign sin[228]  =  8'b11000001;     //228pi/512
  assign cos[228]  =  8'b00001010;     //228pi/512
  assign sin[229]  =  8'b11000001;     //229pi/512
  assign cos[229]  =  8'b00001010;     //229pi/512
  assign sin[230]  =  8'b11000001;     //230pi/512
  assign cos[230]  =  8'b00001010;     //230pi/512
  assign sin[231]  =  8'b11000001;     //231pi/512
  assign cos[231]  =  8'b00001001;     //231pi/512
  assign sin[232]  =  8'b11000001;     //232pi/512
  assign cos[232]  =  8'b00001001;     //232pi/512
  assign sin[233]  =  8'b11000001;     //233pi/512
  assign cos[233]  =  8'b00001001;     //233pi/512
  assign sin[234]  =  8'b11000001;     //234pi/512
  assign cos[234]  =  8'b00001000;     //234pi/512
  assign sin[235]  =  8'b11000001;     //235pi/512
  assign cos[235]  =  8'b00001000;     //235pi/512
  assign sin[236]  =  8'b11000000;     //236pi/512
  assign cos[236]  =  8'b00000111;     //236pi/512
  assign sin[237]  =  8'b11000000;     //237pi/512
  assign cos[237]  =  8'b00000111;     //237pi/512
  assign sin[238]  =  8'b11000000;     //238pi/512
  assign cos[238]  =  8'b00000111;     //238pi/512
  assign sin[239]  =  8'b11000000;     //239pi/512
  assign cos[239]  =  8'b00000110;     //239pi/512
  assign sin[240]  =  8'b11000000;     //240pi/512
  assign cos[240]  =  8'b00000110;     //240pi/512
  assign sin[241]  =  8'b11000000;     //241pi/512
  assign cos[241]  =  8'b00000101;     //241pi/512
  assign sin[242]  =  8'b11000000;     //242pi/512
  assign cos[242]  =  8'b00000101;     //242pi/512
  assign sin[243]  =  8'b11000000;     //243pi/512
  assign cos[243]  =  8'b00000101;     //243pi/512
  assign sin[244]  =  8'b11000000;     //244pi/512
  assign cos[244]  =  8'b00000100;     //244pi/512
  assign sin[245]  =  8'b11000000;     //245pi/512
  assign cos[245]  =  8'b00000100;     //245pi/512
  assign sin[246]  =  8'b11000000;     //246pi/512
  assign cos[246]  =  8'b00000011;     //246pi/512
  assign sin[247]  =  8'b11000000;     //247pi/512
  assign cos[247]  =  8'b00000011;     //247pi/512
  assign sin[248]  =  8'b11000000;     //248pi/512
  assign cos[248]  =  8'b00000011;     //248pi/512
  assign sin[249]  =  8'b11000000;     //249pi/512
  assign cos[249]  =  8'b00000010;     //249pi/512
  assign sin[250]  =  8'b11000000;     //250pi/512
  assign cos[250]  =  8'b00000010;     //250pi/512
  assign sin[251]  =  8'b11000000;     //251pi/512
  assign cos[251]  =  8'b00000001;     //251pi/512
  assign sin[252]  =  8'b11000000;     //252pi/512
  assign cos[252]  =  8'b00000001;     //252pi/512
  assign sin[253]  =  8'b11000000;     //253pi/512
  assign cos[253]  =  8'b00000001;     //253pi/512
  assign sin[254]  =  8'b11000000;     //254pi/512
  assign cos[254]  =  8'b00000000;     //254pi/512
  assign sin[255]  =  8'b11000000;     //255pi/512
  assign cos[255]  =  8'b00000000;     //255pi/512
  assign sin[256]  =  8'b11000000;     //256pi/512
  assign cos[256]  =  8'b00000000;     //256pi/512
  assign sin[257]  =  8'b11000000;     //257pi/512
  assign cos[257]  =  8'b00000000;     //257pi/512
  assign sin[258]  =  8'b11000000;     //258pi/512
  assign cos[258]  =  8'b11111111;     //258pi/512
  assign sin[259]  =  8'b11000000;     //259pi/512
  assign cos[259]  =  8'b11111111;     //259pi/512
  assign sin[260]  =  8'b11000000;     //260pi/512
  assign cos[260]  =  8'b11111110;     //260pi/512
  assign sin[261]  =  8'b11000000;     //261pi/512
  assign cos[261]  =  8'b11111110;     //261pi/512
  assign sin[262]  =  8'b11000000;     //262pi/512
  assign cos[262]  =  8'b11111110;     //262pi/512
  assign sin[263]  =  8'b11000000;     //263pi/512
  assign cos[263]  =  8'b11111101;     //263pi/512
  assign sin[264]  =  8'b11000000;     //264pi/512
  assign cos[264]  =  8'b11111101;     //264pi/512
  assign sin[265]  =  8'b11000000;     //265pi/512
  assign cos[265]  =  8'b11111100;     //265pi/512
  assign sin[266]  =  8'b11000000;     //266pi/512
  assign cos[266]  =  8'b11111100;     //266pi/512
  assign sin[267]  =  8'b11000000;     //267pi/512
  assign cos[267]  =  8'b11111100;     //267pi/512
  assign sin[268]  =  8'b11000000;     //268pi/512
  assign cos[268]  =  8'b11111011;     //268pi/512
  assign sin[269]  =  8'b11000000;     //269pi/512
  assign cos[269]  =  8'b11111011;     //269pi/512
  assign sin[270]  =  8'b11000000;     //270pi/512
  assign cos[270]  =  8'b11111011;     //270pi/512
  assign sin[271]  =  8'b11000000;     //271pi/512
  assign cos[271]  =  8'b11111010;     //271pi/512
  assign sin[272]  =  8'b11000000;     //272pi/512
  assign cos[272]  =  8'b11111010;     //272pi/512
  assign sin[273]  =  8'b11000000;     //273pi/512
  assign cos[273]  =  8'b11111001;     //273pi/512
  assign sin[274]  =  8'b11000000;     //274pi/512
  assign cos[274]  =  8'b11111001;     //274pi/512
  assign sin[275]  =  8'b11000000;     //275pi/512
  assign cos[275]  =  8'b11111001;     //275pi/512
  assign sin[276]  =  8'b11000000;     //276pi/512
  assign cos[276]  =  8'b11111000;     //276pi/512
  assign sin[277]  =  8'b11000001;     //277pi/512
  assign cos[277]  =  8'b11111000;     //277pi/512
  assign sin[278]  =  8'b11000001;     //278pi/512
  assign cos[278]  =  8'b11110111;     //278pi/512
  assign sin[279]  =  8'b11000001;     //279pi/512
  assign cos[279]  =  8'b11110111;     //279pi/512
  assign sin[280]  =  8'b11000001;     //280pi/512
  assign cos[280]  =  8'b11110111;     //280pi/512
  assign sin[281]  =  8'b11000001;     //281pi/512
  assign cos[281]  =  8'b11110110;     //281pi/512
  assign sin[282]  =  8'b11000001;     //282pi/512
  assign cos[282]  =  8'b11110110;     //282pi/512
  assign sin[283]  =  8'b11000001;     //283pi/512
  assign cos[283]  =  8'b11110101;     //283pi/512
  assign sin[284]  =  8'b11000001;     //284pi/512
  assign cos[284]  =  8'b11110101;     //284pi/512
  assign sin[285]  =  8'b11000001;     //285pi/512
  assign cos[285]  =  8'b11110101;     //285pi/512
  assign sin[286]  =  8'b11000001;     //286pi/512
  assign cos[286]  =  8'b11110100;     //286pi/512
  assign sin[287]  =  8'b11000001;     //287pi/512
  assign cos[287]  =  8'b11110100;     //287pi/512
  assign sin[288]  =  8'b11000001;     //288pi/512
  assign cos[288]  =  8'b11110100;     //288pi/512
  assign sin[289]  =  8'b11000001;     //289pi/512
  assign cos[289]  =  8'b11110011;     //289pi/512
  assign sin[290]  =  8'b11000001;     //290pi/512
  assign cos[290]  =  8'b11110011;     //290pi/512
  assign sin[291]  =  8'b11000001;     //291pi/512
  assign cos[291]  =  8'b11110010;     //291pi/512
  assign sin[292]  =  8'b11000010;     //292pi/512
  assign cos[292]  =  8'b11110010;     //292pi/512
  assign sin[293]  =  8'b11000010;     //293pi/512
  assign cos[293]  =  8'b11110010;     //293pi/512
  assign sin[294]  =  8'b11000010;     //294pi/512
  assign cos[294]  =  8'b11110001;     //294pi/512
  assign sin[295]  =  8'b11000010;     //295pi/512
  assign cos[295]  =  8'b11110001;     //295pi/512
  assign sin[296]  =  8'b11000010;     //296pi/512
  assign cos[296]  =  8'b11110000;     //296pi/512
  assign sin[297]  =  8'b11000010;     //297pi/512
  assign cos[297]  =  8'b11110000;     //297pi/512
  assign sin[298]  =  8'b11000010;     //298pi/512
  assign cos[298]  =  8'b11110000;     //298pi/512
  assign sin[299]  =  8'b11000010;     //299pi/512
  assign cos[299]  =  8'b11101111;     //299pi/512
  assign sin[300]  =  8'b11000010;     //300pi/512
  assign cos[300]  =  8'b11101111;     //300pi/512
  assign sin[301]  =  8'b11000010;     //301pi/512
  assign cos[301]  =  8'b11101111;     //301pi/512
  assign sin[302]  =  8'b11000011;     //302pi/512
  assign cos[302]  =  8'b11101110;     //302pi/512
  assign sin[303]  =  8'b11000011;     //303pi/512
  assign cos[303]  =  8'b11101110;     //303pi/512
  assign sin[304]  =  8'b11000011;     //304pi/512
  assign cos[304]  =  8'b11101101;     //304pi/512
  assign sin[305]  =  8'b11000011;     //305pi/512
  assign cos[305]  =  8'b11101101;     //305pi/512
  assign sin[306]  =  8'b11000011;     //306pi/512
  assign cos[306]  =  8'b11101101;     //306pi/512
  assign sin[307]  =  8'b11000011;     //307pi/512
  assign cos[307]  =  8'b11101100;     //307pi/512
  assign sin[308]  =  8'b11000011;     //308pi/512
  assign cos[308]  =  8'b11101100;     //308pi/512
  assign sin[309]  =  8'b11000011;     //309pi/512
  assign cos[309]  =  8'b11101100;     //309pi/512
  assign sin[310]  =  8'b11000011;     //310pi/512
  assign cos[310]  =  8'b11101011;     //310pi/512
  assign sin[311]  =  8'b11000100;     //311pi/512
  assign cos[311]  =  8'b11101011;     //311pi/512
  assign sin[312]  =  8'b11000100;     //312pi/512
  assign cos[312]  =  8'b11101010;     //312pi/512
  assign sin[313]  =  8'b11000100;     //313pi/512
  assign cos[313]  =  8'b11101010;     //313pi/512
  assign sin[314]  =  8'b11000100;     //314pi/512
  assign cos[314]  =  8'b11101010;     //314pi/512
  assign sin[315]  =  8'b11000100;     //315pi/512
  assign cos[315]  =  8'b11101001;     //315pi/512
  assign sin[316]  =  8'b11000100;     //316pi/512
  assign cos[316]  =  8'b11101001;     //316pi/512
  assign sin[317]  =  8'b11000100;     //317pi/512
  assign cos[317]  =  8'b11101001;     //317pi/512
  assign sin[318]  =  8'b11000101;     //318pi/512
  assign cos[318]  =  8'b11101000;     //318pi/512
  assign sin[319]  =  8'b11000101;     //319pi/512
  assign cos[319]  =  8'b11101000;     //319pi/512
  assign sin[320]  =  8'b11000101;     //320pi/512
  assign cos[320]  =  8'b11101000;     //320pi/512
  assign sin[321]  =  8'b11000101;     //321pi/512
  assign cos[321]  =  8'b11100111;     //321pi/512
  assign sin[322]  =  8'b11000101;     //322pi/512
  assign cos[322]  =  8'b11100111;     //322pi/512
  assign sin[323]  =  8'b11000101;     //323pi/512
  assign cos[323]  =  8'b11100110;     //323pi/512
  assign sin[324]  =  8'b11000101;     //324pi/512
  assign cos[324]  =  8'b11100110;     //324pi/512
  assign sin[325]  =  8'b11000110;     //325pi/512
  assign cos[325]  =  8'b11100110;     //325pi/512
  assign sin[326]  =  8'b11000110;     //326pi/512
  assign cos[326]  =  8'b11100101;     //326pi/512
  assign sin[327]  =  8'b11000110;     //327pi/512
  assign cos[327]  =  8'b11100101;     //327pi/512
  assign sin[328]  =  8'b11000110;     //328pi/512
  assign cos[328]  =  8'b11100101;     //328pi/512
  assign sin[329]  =  8'b11000110;     //329pi/512
  assign cos[329]  =  8'b11100100;     //329pi/512
  assign sin[330]  =  8'b11000110;     //330pi/512
  assign cos[330]  =  8'b11100100;     //330pi/512
  assign sin[331]  =  8'b11000111;     //331pi/512
  assign cos[331]  =  8'b11100100;     //331pi/512
  assign sin[332]  =  8'b11000111;     //332pi/512
  assign cos[332]  =  8'b11100011;     //332pi/512
  assign sin[333]  =  8'b11000111;     //333pi/512
  assign cos[333]  =  8'b11100011;     //333pi/512
  assign sin[334]  =  8'b11000111;     //334pi/512
  assign cos[334]  =  8'b11100011;     //334pi/512
  assign sin[335]  =  8'b11000111;     //335pi/512
  assign cos[335]  =  8'b11100010;     //335pi/512
  assign sin[336]  =  8'b11001000;     //336pi/512
  assign cos[336]  =  8'b11100010;     //336pi/512
  assign sin[337]  =  8'b11001000;     //337pi/512
  assign cos[337]  =  8'b11100001;     //337pi/512
  assign sin[338]  =  8'b11001000;     //338pi/512
  assign cos[338]  =  8'b11100001;     //338pi/512
  assign sin[339]  =  8'b11001000;     //339pi/512
  assign cos[339]  =  8'b11100001;     //339pi/512
  assign sin[340]  =  8'b11001000;     //340pi/512
  assign cos[340]  =  8'b11100000;     //340pi/512
  assign sin[341]  =  8'b11001001;     //341pi/512
  assign cos[341]  =  8'b11100000;     //341pi/512
  assign sin[342]  =  8'b11001001;     //342pi/512
  assign cos[342]  =  8'b11100000;     //342pi/512
  assign sin[343]  =  8'b11001001;     //343pi/512
  assign cos[343]  =  8'b11011111;     //343pi/512
  assign sin[344]  =  8'b11001001;     //344pi/512
  assign cos[344]  =  8'b11011111;     //344pi/512
  assign sin[345]  =  8'b11001001;     //345pi/512
  assign cos[345]  =  8'b11011111;     //345pi/512
  assign sin[346]  =  8'b11001010;     //346pi/512
  assign cos[346]  =  8'b11011110;     //346pi/512
  assign sin[347]  =  8'b11001010;     //347pi/512
  assign cos[347]  =  8'b11011110;     //347pi/512
  assign sin[348]  =  8'b11001010;     //348pi/512
  assign cos[348]  =  8'b11011110;     //348pi/512
  assign sin[349]  =  8'b11001010;     //349pi/512
  assign cos[349]  =  8'b11011101;     //349pi/512
  assign sin[350]  =  8'b11001010;     //350pi/512
  assign cos[350]  =  8'b11011101;     //350pi/512
  assign sin[351]  =  8'b11001011;     //351pi/512
  assign cos[351]  =  8'b11011101;     //351pi/512
  assign sin[352]  =  8'b11001011;     //352pi/512
  assign cos[352]  =  8'b11011100;     //352pi/512
  assign sin[353]  =  8'b11001011;     //353pi/512
  assign cos[353]  =  8'b11011100;     //353pi/512
  assign sin[354]  =  8'b11001011;     //354pi/512
  assign cos[354]  =  8'b11011100;     //354pi/512
  assign sin[355]  =  8'b11001011;     //355pi/512
  assign cos[355]  =  8'b11011011;     //355pi/512
  assign sin[356]  =  8'b11001100;     //356pi/512
  assign cos[356]  =  8'b11011011;     //356pi/512
  assign sin[357]  =  8'b11001100;     //357pi/512
  assign cos[357]  =  8'b11011011;     //357pi/512
  assign sin[358]  =  8'b11001100;     //358pi/512
  assign cos[358]  =  8'b11011011;     //358pi/512
  assign sin[359]  =  8'b11001100;     //359pi/512
  assign cos[359]  =  8'b11011010;     //359pi/512
  assign sin[360]  =  8'b11001101;     //360pi/512
  assign cos[360]  =  8'b11011010;     //360pi/512
  assign sin[361]  =  8'b11001101;     //361pi/512
  assign cos[361]  =  8'b11011010;     //361pi/512
  assign sin[362]  =  8'b11001101;     //362pi/512
  assign cos[362]  =  8'b11011001;     //362pi/512
  assign sin[363]  =  8'b11001101;     //363pi/512
  assign cos[363]  =  8'b11011001;     //363pi/512
  assign sin[364]  =  8'b11001110;     //364pi/512
  assign cos[364]  =  8'b11011001;     //364pi/512
  assign sin[365]  =  8'b11001110;     //365pi/512
  assign cos[365]  =  8'b11011000;     //365pi/512
  assign sin[366]  =  8'b11001110;     //366pi/512
  assign cos[366]  =  8'b11011000;     //366pi/512
  assign sin[367]  =  8'b11001110;     //367pi/512
  assign cos[367]  =  8'b11011000;     //367pi/512
  assign sin[368]  =  8'b11001111;     //368pi/512
  assign cos[368]  =  8'b11010111;     //368pi/512
  assign sin[369]  =  8'b11001111;     //369pi/512
  assign cos[369]  =  8'b11010111;     //369pi/512
  assign sin[370]  =  8'b11001111;     //370pi/512
  assign cos[370]  =  8'b11010111;     //370pi/512
  assign sin[371]  =  8'b11001111;     //371pi/512
  assign cos[371]  =  8'b11010110;     //371pi/512
  assign sin[372]  =  8'b11010000;     //372pi/512
  assign cos[372]  =  8'b11010110;     //372pi/512
  assign sin[373]  =  8'b11010000;     //373pi/512
  assign cos[373]  =  8'b11010110;     //373pi/512
  assign sin[374]  =  8'b11010000;     //374pi/512
  assign cos[374]  =  8'b11010110;     //374pi/512
  assign sin[375]  =  8'b11010000;     //375pi/512
  assign cos[375]  =  8'b11010101;     //375pi/512
  assign sin[376]  =  8'b11010001;     //376pi/512
  assign cos[376]  =  8'b11010101;     //376pi/512
  assign sin[377]  =  8'b11010001;     //377pi/512
  assign cos[377]  =  8'b11010101;     //377pi/512
  assign sin[378]  =  8'b11010001;     //378pi/512
  assign cos[378]  =  8'b11010100;     //378pi/512
  assign sin[379]  =  8'b11010001;     //379pi/512
  assign cos[379]  =  8'b11010100;     //379pi/512
  assign sin[380]  =  8'b11010010;     //380pi/512
  assign cos[380]  =  8'b11010100;     //380pi/512
  assign sin[381]  =  8'b11010010;     //381pi/512
  assign cos[381]  =  8'b11010100;     //381pi/512
  assign sin[382]  =  8'b11010010;     //382pi/512
  assign cos[382]  =  8'b11010011;     //382pi/512
  assign sin[383]  =  8'b11010010;     //383pi/512
  assign cos[383]  =  8'b11010011;     //383pi/512
  assign sin[384]  =  8'b11010011;     //384pi/512
  assign cos[384]  =  8'b11010011;     //384pi/512
  assign sin[385]  =  8'b11010011;     //385pi/512
  assign cos[385]  =  8'b11010010;     //385pi/512
  assign sin[386]  =  8'b11010011;     //386pi/512
  assign cos[386]  =  8'b11010010;     //386pi/512
  assign sin[387]  =  8'b11010100;     //387pi/512
  assign cos[387]  =  8'b11010010;     //387pi/512
  assign sin[388]  =  8'b11010100;     //388pi/512
  assign cos[388]  =  8'b11010010;     //388pi/512
  assign sin[389]  =  8'b11010100;     //389pi/512
  assign cos[389]  =  8'b11010001;     //389pi/512
  assign sin[390]  =  8'b11010100;     //390pi/512
  assign cos[390]  =  8'b11010001;     //390pi/512
  assign sin[391]  =  8'b11010101;     //391pi/512
  assign cos[391]  =  8'b11010001;     //391pi/512
  assign sin[392]  =  8'b11010101;     //392pi/512
  assign cos[392]  =  8'b11010001;     //392pi/512
  assign sin[393]  =  8'b11010101;     //393pi/512
  assign cos[393]  =  8'b11010000;     //393pi/512
  assign sin[394]  =  8'b11010110;     //394pi/512
  assign cos[394]  =  8'b11010000;     //394pi/512
  assign sin[395]  =  8'b11010110;     //395pi/512
  assign cos[395]  =  8'b11010000;     //395pi/512
  assign sin[396]  =  8'b11010110;     //396pi/512
  assign cos[396]  =  8'b11010000;     //396pi/512
  assign sin[397]  =  8'b11010110;     //397pi/512
  assign cos[397]  =  8'b11001111;     //397pi/512
  assign sin[398]  =  8'b11010111;     //398pi/512
  assign cos[398]  =  8'b11001111;     //398pi/512
  assign sin[399]  =  8'b11010111;     //399pi/512
  assign cos[399]  =  8'b11001111;     //399pi/512
  assign sin[400]  =  8'b11010111;     //400pi/512
  assign cos[400]  =  8'b11001111;     //400pi/512
  assign sin[401]  =  8'b11011000;     //401pi/512
  assign cos[401]  =  8'b11001110;     //401pi/512
  assign sin[402]  =  8'b11011000;     //402pi/512
  assign cos[402]  =  8'b11001110;     //402pi/512
  assign sin[403]  =  8'b11011000;     //403pi/512
  assign cos[403]  =  8'b11001110;     //403pi/512
  assign sin[404]  =  8'b11011001;     //404pi/512
  assign cos[404]  =  8'b11001110;     //404pi/512
  assign sin[405]  =  8'b11011001;     //405pi/512
  assign cos[405]  =  8'b11001101;     //405pi/512
  assign sin[406]  =  8'b11011001;     //406pi/512
  assign cos[406]  =  8'b11001101;     //406pi/512
  assign sin[407]  =  8'b11011010;     //407pi/512
  assign cos[407]  =  8'b11001101;     //407pi/512
  assign sin[408]  =  8'b11011010;     //408pi/512
  assign cos[408]  =  8'b11001101;     //408pi/512
  assign sin[409]  =  8'b11011010;     //409pi/512
  assign cos[409]  =  8'b11001100;     //409pi/512
  assign sin[410]  =  8'b11011011;     //410pi/512
  assign cos[410]  =  8'b11001100;     //410pi/512
  assign sin[411]  =  8'b11011011;     //411pi/512
  assign cos[411]  =  8'b11001100;     //411pi/512
  assign sin[412]  =  8'b11011011;     //412pi/512
  assign cos[412]  =  8'b11001100;     //412pi/512
  assign sin[413]  =  8'b11011011;     //413pi/512
  assign cos[413]  =  8'b11001011;     //413pi/512
  assign sin[414]  =  8'b11011100;     //414pi/512
  assign cos[414]  =  8'b11001011;     //414pi/512
  assign sin[415]  =  8'b11011100;     //415pi/512
  assign cos[415]  =  8'b11001011;     //415pi/512
  assign sin[416]  =  8'b11011100;     //416pi/512
  assign cos[416]  =  8'b11001011;     //416pi/512
  assign sin[417]  =  8'b11011101;     //417pi/512
  assign cos[417]  =  8'b11001011;     //417pi/512
  assign sin[418]  =  8'b11011101;     //418pi/512
  assign cos[418]  =  8'b11001010;     //418pi/512
  assign sin[419]  =  8'b11011101;     //419pi/512
  assign cos[419]  =  8'b11001010;     //419pi/512
  assign sin[420]  =  8'b11011110;     //420pi/512
  assign cos[420]  =  8'b11001010;     //420pi/512
  assign sin[421]  =  8'b11011110;     //421pi/512
  assign cos[421]  =  8'b11001010;     //421pi/512
  assign sin[422]  =  8'b11011110;     //422pi/512
  assign cos[422]  =  8'b11001010;     //422pi/512
  assign sin[423]  =  8'b11011111;     //423pi/512
  assign cos[423]  =  8'b11001001;     //423pi/512
  assign sin[424]  =  8'b11011111;     //424pi/512
  assign cos[424]  =  8'b11001001;     //424pi/512
  assign sin[425]  =  8'b11011111;     //425pi/512
  assign cos[425]  =  8'b11001001;     //425pi/512
  assign sin[426]  =  8'b11100000;     //426pi/512
  assign cos[426]  =  8'b11001001;     //426pi/512
  assign sin[427]  =  8'b11100000;     //427pi/512
  assign cos[427]  =  8'b11001001;     //427pi/512
  assign sin[428]  =  8'b11100000;     //428pi/512
  assign cos[428]  =  8'b11001000;     //428pi/512
  assign sin[429]  =  8'b11100001;     //429pi/512
  assign cos[429]  =  8'b11001000;     //429pi/512
  assign sin[430]  =  8'b11100001;     //430pi/512
  assign cos[430]  =  8'b11001000;     //430pi/512
  assign sin[431]  =  8'b11100001;     //431pi/512
  assign cos[431]  =  8'b11001000;     //431pi/512
  assign sin[432]  =  8'b11100010;     //432pi/512
  assign cos[432]  =  8'b11001000;     //432pi/512
  assign sin[433]  =  8'b11100010;     //433pi/512
  assign cos[433]  =  8'b11000111;     //433pi/512
  assign sin[434]  =  8'b11100011;     //434pi/512
  assign cos[434]  =  8'b11000111;     //434pi/512
  assign sin[435]  =  8'b11100011;     //435pi/512
  assign cos[435]  =  8'b11000111;     //435pi/512
  assign sin[436]  =  8'b11100011;     //436pi/512
  assign cos[436]  =  8'b11000111;     //436pi/512
  assign sin[437]  =  8'b11100100;     //437pi/512
  assign cos[437]  =  8'b11000111;     //437pi/512
  assign sin[438]  =  8'b11100100;     //438pi/512
  assign cos[438]  =  8'b11000110;     //438pi/512
  assign sin[439]  =  8'b11100100;     //439pi/512
  assign cos[439]  =  8'b11000110;     //439pi/512
  assign sin[440]  =  8'b11100101;     //440pi/512
  assign cos[440]  =  8'b11000110;     //440pi/512
  assign sin[441]  =  8'b11100101;     //441pi/512
  assign cos[441]  =  8'b11000110;     //441pi/512
  assign sin[442]  =  8'b11100101;     //442pi/512
  assign cos[442]  =  8'b11000110;     //442pi/512
  assign sin[443]  =  8'b11100110;     //443pi/512
  assign cos[443]  =  8'b11000110;     //443pi/512
  assign sin[444]  =  8'b11100110;     //444pi/512
  assign cos[444]  =  8'b11000101;     //444pi/512
  assign sin[445]  =  8'b11100110;     //445pi/512
  assign cos[445]  =  8'b11000101;     //445pi/512
  assign sin[446]  =  8'b11100111;     //446pi/512
  assign cos[446]  =  8'b11000101;     //446pi/512
  assign sin[447]  =  8'b11100111;     //447pi/512
  assign cos[447]  =  8'b11000101;     //447pi/512
  assign sin[448]  =  8'b11101000;     //448pi/512
  assign cos[448]  =  8'b11000101;     //448pi/512
  assign sin[449]  =  8'b11101000;     //449pi/512
  assign cos[449]  =  8'b11000101;     //449pi/512
  assign sin[450]  =  8'b11101000;     //450pi/512
  assign cos[450]  =  8'b11000101;     //450pi/512
  assign sin[451]  =  8'b11101001;     //451pi/512
  assign cos[451]  =  8'b11000100;     //451pi/512
  assign sin[452]  =  8'b11101001;     //452pi/512
  assign cos[452]  =  8'b11000100;     //452pi/512
  assign sin[453]  =  8'b11101001;     //453pi/512
  assign cos[453]  =  8'b11000100;     //453pi/512
  assign sin[454]  =  8'b11101010;     //454pi/512
  assign cos[454]  =  8'b11000100;     //454pi/512
  assign sin[455]  =  8'b11101010;     //455pi/512
  assign cos[455]  =  8'b11000100;     //455pi/512
  assign sin[456]  =  8'b11101010;     //456pi/512
  assign cos[456]  =  8'b11000100;     //456pi/512
  assign sin[457]  =  8'b11101011;     //457pi/512
  assign cos[457]  =  8'b11000100;     //457pi/512
  assign sin[458]  =  8'b11101011;     //458pi/512
  assign cos[458]  =  8'b11000011;     //458pi/512
  assign sin[459]  =  8'b11101100;     //459pi/512
  assign cos[459]  =  8'b11000011;     //459pi/512
  assign sin[460]  =  8'b11101100;     //460pi/512
  assign cos[460]  =  8'b11000011;     //460pi/512
  assign sin[461]  =  8'b11101100;     //461pi/512
  assign cos[461]  =  8'b11000011;     //461pi/512
  assign sin[462]  =  8'b11101101;     //462pi/512
  assign cos[462]  =  8'b11000011;     //462pi/512
  assign sin[463]  =  8'b11101101;     //463pi/512
  assign cos[463]  =  8'b11000011;     //463pi/512
  assign sin[464]  =  8'b11101101;     //464pi/512
  assign cos[464]  =  8'b11000011;     //464pi/512
  assign sin[465]  =  8'b11101110;     //465pi/512
  assign cos[465]  =  8'b11000011;     //465pi/512
  assign sin[466]  =  8'b11101110;     //466pi/512
  assign cos[466]  =  8'b11000011;     //466pi/512
  assign sin[467]  =  8'b11101111;     //467pi/512
  assign cos[467]  =  8'b11000010;     //467pi/512
  assign sin[468]  =  8'b11101111;     //468pi/512
  assign cos[468]  =  8'b11000010;     //468pi/512
  assign sin[469]  =  8'b11101111;     //469pi/512
  assign cos[469]  =  8'b11000010;     //469pi/512
  assign sin[470]  =  8'b11110000;     //470pi/512
  assign cos[470]  =  8'b11000010;     //470pi/512
  assign sin[471]  =  8'b11110000;     //471pi/512
  assign cos[471]  =  8'b11000010;     //471pi/512
  assign sin[472]  =  8'b11110000;     //472pi/512
  assign cos[472]  =  8'b11000010;     //472pi/512
  assign sin[473]  =  8'b11110001;     //473pi/512
  assign cos[473]  =  8'b11000010;     //473pi/512
  assign sin[474]  =  8'b11110001;     //474pi/512
  assign cos[474]  =  8'b11000010;     //474pi/512
  assign sin[475]  =  8'b11110010;     //475pi/512
  assign cos[475]  =  8'b11000010;     //475pi/512
  assign sin[476]  =  8'b11110010;     //476pi/512
  assign cos[476]  =  8'b11000010;     //476pi/512
  assign sin[477]  =  8'b11110010;     //477pi/512
  assign cos[477]  =  8'b11000001;     //477pi/512
  assign sin[478]  =  8'b11110011;     //478pi/512
  assign cos[478]  =  8'b11000001;     //478pi/512
  assign sin[479]  =  8'b11110011;     //479pi/512
  assign cos[479]  =  8'b11000001;     //479pi/512
  assign sin[480]  =  8'b11110100;     //480pi/512
  assign cos[480]  =  8'b11000001;     //480pi/512
  assign sin[481]  =  8'b11110100;     //481pi/512
  assign cos[481]  =  8'b11000001;     //481pi/512
  assign sin[482]  =  8'b11110100;     //482pi/512
  assign cos[482]  =  8'b11000001;     //482pi/512
  assign sin[483]  =  8'b11110101;     //483pi/512
  assign cos[483]  =  8'b11000001;     //483pi/512
  assign sin[484]  =  8'b11110101;     //484pi/512
  assign cos[484]  =  8'b11000001;     //484pi/512
  assign sin[485]  =  8'b11110101;     //485pi/512
  assign cos[485]  =  8'b11000001;     //485pi/512
  assign sin[486]  =  8'b11110110;     //486pi/512
  assign cos[486]  =  8'b11000001;     //486pi/512
  assign sin[487]  =  8'b11110110;     //487pi/512
  assign cos[487]  =  8'b11000001;     //487pi/512
  assign sin[488]  =  8'b11110111;     //488pi/512
  assign cos[488]  =  8'b11000001;     //488pi/512
  assign sin[489]  =  8'b11110111;     //489pi/512
  assign cos[489]  =  8'b11000001;     //489pi/512
  assign sin[490]  =  8'b11110111;     //490pi/512
  assign cos[490]  =  8'b11000001;     //490pi/512
  assign sin[491]  =  8'b11111000;     //491pi/512
  assign cos[491]  =  8'b11000001;     //491pi/512
  assign sin[492]  =  8'b11111000;     //492pi/512
  assign cos[492]  =  8'b11000000;     //492pi/512
  assign sin[493]  =  8'b11111001;     //493pi/512
  assign cos[493]  =  8'b11000000;     //493pi/512
  assign sin[494]  =  8'b11111001;     //494pi/512
  assign cos[494]  =  8'b11000000;     //494pi/512
  assign sin[495]  =  8'b11111001;     //495pi/512
  assign cos[495]  =  8'b11000000;     //495pi/512
  assign sin[496]  =  8'b11111010;     //496pi/512
  assign cos[496]  =  8'b11000000;     //496pi/512
  assign sin[497]  =  8'b11111010;     //497pi/512
  assign cos[497]  =  8'b11000000;     //497pi/512
  assign sin[498]  =  8'b11111011;     //498pi/512
  assign cos[498]  =  8'b11000000;     //498pi/512
  assign sin[499]  =  8'b11111011;     //499pi/512
  assign cos[499]  =  8'b11000000;     //499pi/512
  assign sin[500]  =  8'b11111011;     //500pi/512
  assign cos[500]  =  8'b11000000;     //500pi/512
  assign sin[501]  =  8'b11111100;     //501pi/512
  assign cos[501]  =  8'b11000000;     //501pi/512
  assign sin[502]  =  8'b11111100;     //502pi/512
  assign cos[502]  =  8'b11000000;     //502pi/512
  assign sin[503]  =  8'b11111100;     //503pi/512
  assign cos[503]  =  8'b11000000;     //503pi/512
  assign sin[504]  =  8'b11111101;     //504pi/512
  assign cos[504]  =  8'b11000000;     //504pi/512
  assign sin[505]  =  8'b11111101;     //505pi/512
  assign cos[505]  =  8'b11000000;     //505pi/512
  assign sin[506]  =  8'b11111110;     //506pi/512
  assign cos[506]  =  8'b11000000;     //506pi/512
  assign sin[507]  =  8'b11111110;     //507pi/512
  assign cos[507]  =  8'b11000000;     //507pi/512
  assign sin[508]  =  8'b11111110;     //508pi/512
  assign cos[508]  =  8'b11000000;     //508pi/512
  assign sin[509]  =  8'b11111111;     //509pi/512
  assign cos[509]  =  8'b11000000;     //509pi/512
  assign sin[510]  =  8'b11111111;     //510pi/512
  assign cos[510]  =  8'b11000000;     //510pi/512
  assign sin[511]  =  8'b00000000;     //511pi/512
  assign cos[511]  =  8'b11000000;     //511pi/512
/////////////////////////////////////////////////////////////////

  assign sin2[0]  =  8'b00000000;     //0pi/512
  assign cos2[0]  =  8'b01000000;     //0pi/512
  assign sin2[1]  =  8'b00000000;     //1pi/512
  assign cos2[1]  =  8'b00111111;     //1pi/512
  assign sin2[2]  =  8'b11111111;     //2pi/512
  assign cos2[2]  =  8'b00111111;     //2pi/512
  assign sin2[3]  =  8'b11111111;     //3pi/512
  assign cos2[3]  =  8'b00111111;     //3pi/512
  assign sin2[4]  =  8'b11111111;     //4pi/512
  assign cos2[4]  =  8'b00111111;     //4pi/512
  assign sin2[5]  =  8'b11111110;     //5pi/512
  assign cos2[5]  =  8'b00111111;     //5pi/512
  assign sin2[6]  =  8'b11111110;     //6pi/512
  assign cos2[6]  =  8'b00111111;     //6pi/512
  assign sin2[7]  =  8'b11111110;     //7pi/512
  assign cos2[7]  =  8'b00111111;     //7pi/512
  assign sin2[8]  =  8'b11111101;     //8pi/512
  assign cos2[8]  =  8'b00111111;     //8pi/512
  assign sin2[9]  =  8'b11111101;     //9pi/512
  assign cos2[9]  =  8'b00111111;     //9pi/512
  assign sin2[10]  =  8'b11111101;     //10pi/512
  assign cos2[10]  =  8'b00111111;     //10pi/512
  assign sin2[11]  =  8'b11111101;     //11pi/512
  assign cos2[11]  =  8'b00111111;     //11pi/512
  assign sin2[12]  =  8'b11111100;     //12pi/512
  assign cos2[12]  =  8'b00111111;     //12pi/512
  assign sin2[13]  =  8'b11111100;     //13pi/512
  assign cos2[13]  =  8'b00111111;     //13pi/512
  assign sin2[14]  =  8'b11111100;     //14pi/512
  assign cos2[14]  =  8'b00111111;     //14pi/512
  assign sin2[15]  =  8'b11111011;     //15pi/512
  assign cos2[15]  =  8'b00111111;     //15pi/512
  assign sin2[16]  =  8'b11111011;     //16pi/512
  assign cos2[16]  =  8'b00111111;     //16pi/512
  assign sin2[17]  =  8'b11111011;     //17pi/512
  assign cos2[17]  =  8'b00111111;     //17pi/512
  assign sin2[18]  =  8'b11111010;     //18pi/512
  assign cos2[18]  =  8'b00111111;     //18pi/512
  assign sin2[19]  =  8'b11111010;     //19pi/512
  assign cos2[19]  =  8'b00111111;     //19pi/512
  assign sin2[20]  =  8'b11111010;     //20pi/512
  assign cos2[20]  =  8'b00111111;     //20pi/512
  assign sin2[21]  =  8'b11111001;     //21pi/512
  assign cos2[21]  =  8'b00111111;     //21pi/512
  assign sin2[22]  =  8'b11111001;     //22pi/512
  assign cos2[22]  =  8'b00111111;     //22pi/512
  assign sin2[23]  =  8'b11111001;     //23pi/512
  assign cos2[23]  =  8'b00111111;     //23pi/512
  assign sin2[24]  =  8'b11111000;     //24pi/512
  assign cos2[24]  =  8'b00111111;     //24pi/512
  assign sin2[25]  =  8'b11111000;     //25pi/512
  assign cos2[25]  =  8'b00111111;     //25pi/512
  assign sin2[26]  =  8'b11111000;     //26pi/512
  assign cos2[26]  =  8'b00111111;     //26pi/512
  assign sin2[27]  =  8'b11111000;     //27pi/512
  assign cos2[27]  =  8'b00111111;     //27pi/512
  assign sin2[28]  =  8'b11110111;     //28pi/512
  assign cos2[28]  =  8'b00111111;     //28pi/512
  assign sin2[29]  =  8'b11110111;     //29pi/512
  assign cos2[29]  =  8'b00111111;     //29pi/512
  assign sin2[30]  =  8'b11110111;     //30pi/512
  assign cos2[30]  =  8'b00111111;     //30pi/512
  assign sin2[31]  =  8'b11110110;     //31pi/512
  assign cos2[31]  =  8'b00111111;     //31pi/512
  assign sin2[32]  =  8'b11110110;     //32pi/512
  assign cos2[32]  =  8'b00111111;     //32pi/512
  assign sin2[33]  =  8'b11110110;     //33pi/512
  assign cos2[33]  =  8'b00111111;     //33pi/512
  assign sin2[34]  =  8'b11110101;     //34pi/512
  assign cos2[34]  =  8'b00111111;     //34pi/512
  assign sin2[35]  =  8'b11110101;     //35pi/512
  assign cos2[35]  =  8'b00111111;     //35pi/512
  assign sin2[36]  =  8'b11110101;     //36pi/512
  assign cos2[36]  =  8'b00111111;     //36pi/512
  assign sin2[37]  =  8'b11110100;     //37pi/512
  assign cos2[37]  =  8'b00111110;     //37pi/512
  assign sin2[38]  =  8'b11110100;     //38pi/512
  assign cos2[38]  =  8'b00111110;     //38pi/512
  assign sin2[39]  =  8'b11110100;     //39pi/512
  assign cos2[39]  =  8'b00111110;     //39pi/512
  assign sin2[40]  =  8'b11110100;     //40pi/512
  assign cos2[40]  =  8'b00111110;     //40pi/512
  assign sin2[41]  =  8'b11110011;     //41pi/512
  assign cos2[41]  =  8'b00111110;     //41pi/512
  assign sin2[42]  =  8'b11110011;     //42pi/512
  assign cos2[42]  =  8'b00111110;     //42pi/512
  assign sin2[43]  =  8'b11110011;     //43pi/512
  assign cos2[43]  =  8'b00111110;     //43pi/512
  assign sin2[44]  =  8'b11110010;     //44pi/512
  assign cos2[44]  =  8'b00111110;     //44pi/512
  assign sin2[45]  =  8'b11110010;     //45pi/512
  assign cos2[45]  =  8'b00111110;     //45pi/512
  assign sin2[46]  =  8'b11110010;     //46pi/512
  assign cos2[46]  =  8'b00111110;     //46pi/512
  assign sin2[47]  =  8'b11110001;     //47pi/512
  assign cos2[47]  =  8'b00111110;     //47pi/512
  assign sin2[48]  =  8'b11110001;     //48pi/512
  assign cos2[48]  =  8'b00111110;     //48pi/512
  assign sin2[49]  =  8'b11110001;     //49pi/512
  assign cos2[49]  =  8'b00111110;     //49pi/512
  assign sin2[50]  =  8'b11110000;     //50pi/512
  assign cos2[50]  =  8'b00111110;     //50pi/512
  assign sin2[51]  =  8'b11110000;     //51pi/512
  assign cos2[51]  =  8'b00111110;     //51pi/512
  assign sin2[52]  =  8'b11110000;     //52pi/512
  assign cos2[52]  =  8'b00111101;     //52pi/512
  assign sin2[53]  =  8'b11110000;     //53pi/512
  assign cos2[53]  =  8'b00111101;     //53pi/512
  assign sin2[54]  =  8'b11101111;     //54pi/512
  assign cos2[54]  =  8'b00111101;     //54pi/512
  assign sin2[55]  =  8'b11101111;     //55pi/512
  assign cos2[55]  =  8'b00111101;     //55pi/512
  assign sin2[56]  =  8'b11101111;     //56pi/512
  assign cos2[56]  =  8'b00111101;     //56pi/512
  assign sin2[57]  =  8'b11101110;     //57pi/512
  assign cos2[57]  =  8'b00111101;     //57pi/512
  assign sin2[58]  =  8'b11101110;     //58pi/512
  assign cos2[58]  =  8'b00111101;     //58pi/512
  assign sin2[59]  =  8'b11101110;     //59pi/512
  assign cos2[59]  =  8'b00111101;     //59pi/512
  assign sin2[60]  =  8'b11101101;     //60pi/512
  assign cos2[60]  =  8'b00111101;     //60pi/512
  assign sin2[61]  =  8'b11101101;     //61pi/512
  assign cos2[61]  =  8'b00111101;     //61pi/512
  assign sin2[62]  =  8'b11101101;     //62pi/512
  assign cos2[62]  =  8'b00111101;     //62pi/512
  assign sin2[63]  =  8'b11101101;     //63pi/512
  assign cos2[63]  =  8'b00111100;     //63pi/512
  assign sin2[64]  =  8'b11101100;     //64pi/512
  assign cos2[64]  =  8'b00111100;     //64pi/512
  assign sin2[65]  =  8'b11101100;     //65pi/512
  assign cos2[65]  =  8'b00111100;     //65pi/512
  assign sin2[66]  =  8'b11101100;     //66pi/512
  assign cos2[66]  =  8'b00111100;     //66pi/512
  assign sin2[67]  =  8'b11101011;     //67pi/512
  assign cos2[67]  =  8'b00111100;     //67pi/512
  assign sin2[68]  =  8'b11101011;     //68pi/512
  assign cos2[68]  =  8'b00111100;     //68pi/512
  assign sin2[69]  =  8'b11101011;     //69pi/512
  assign cos2[69]  =  8'b00111100;     //69pi/512
  assign sin2[70]  =  8'b11101010;     //70pi/512
  assign cos2[70]  =  8'b00111100;     //70pi/512
  assign sin2[71]  =  8'b11101010;     //71pi/512
  assign cos2[71]  =  8'b00111100;     //71pi/512
  assign sin2[72]  =  8'b11101010;     //72pi/512
  assign cos2[72]  =  8'b00111100;     //72pi/512
  assign sin2[73]  =  8'b11101010;     //73pi/512
  assign cos2[73]  =  8'b00111011;     //73pi/512
  assign sin2[74]  =  8'b11101001;     //74pi/512
  assign cos2[74]  =  8'b00111011;     //74pi/512
  assign sin2[75]  =  8'b11101001;     //75pi/512
  assign cos2[75]  =  8'b00111011;     //75pi/512
  assign sin2[76]  =  8'b11101001;     //76pi/512
  assign cos2[76]  =  8'b00111011;     //76pi/512
  assign sin2[77]  =  8'b11101000;     //77pi/512
  assign cos2[77]  =  8'b00111011;     //77pi/512
  assign sin2[78]  =  8'b11101000;     //78pi/512
  assign cos2[78]  =  8'b00111011;     //78pi/512
  assign sin2[79]  =  8'b11101000;     //79pi/512
  assign cos2[79]  =  8'b00111011;     //79pi/512
  assign sin2[80]  =  8'b11101000;     //80pi/512
  assign cos2[80]  =  8'b00111011;     //80pi/512
  assign sin2[81]  =  8'b11100111;     //81pi/512
  assign cos2[81]  =  8'b00111011;     //81pi/512
  assign sin2[82]  =  8'b11100111;     //82pi/512
  assign cos2[82]  =  8'b00111010;     //82pi/512
  assign sin2[83]  =  8'b11100111;     //83pi/512
  assign cos2[83]  =  8'b00111010;     //83pi/512
  assign sin2[84]  =  8'b11100110;     //84pi/512
  assign cos2[84]  =  8'b00111010;     //84pi/512
  assign sin2[85]  =  8'b11100110;     //85pi/512
  assign cos2[85]  =  8'b00111010;     //85pi/512
  assign sin2[86]  =  8'b11100110;     //86pi/512
  assign cos2[86]  =  8'b00111010;     //86pi/512
  assign sin2[87]  =  8'b11100101;     //87pi/512
  assign cos2[87]  =  8'b00111010;     //87pi/512
  assign sin2[88]  =  8'b11100101;     //88pi/512
  assign cos2[88]  =  8'b00111010;     //88pi/512
  assign sin2[89]  =  8'b11100101;     //89pi/512
  assign cos2[89]  =  8'b00111001;     //89pi/512
  assign sin2[90]  =  8'b11100101;     //90pi/512
  assign cos2[90]  =  8'b00111001;     //90pi/512
  assign sin2[91]  =  8'b11100100;     //91pi/512
  assign cos2[91]  =  8'b00111001;     //91pi/512
  assign sin2[92]  =  8'b11100100;     //92pi/512
  assign cos2[92]  =  8'b00111001;     //92pi/512
  assign sin2[93]  =  8'b11100100;     //93pi/512
  assign cos2[93]  =  8'b00111001;     //93pi/512
  assign sin2[94]  =  8'b11100100;     //94pi/512
  assign cos2[94]  =  8'b00111001;     //94pi/512
  assign sin2[95]  =  8'b11100011;     //95pi/512
  assign cos2[95]  =  8'b00111001;     //95pi/512
  assign sin2[96]  =  8'b11100011;     //96pi/512
  assign cos2[96]  =  8'b00111001;     //96pi/512
  assign sin2[97]  =  8'b11100011;     //97pi/512
  assign cos2[97]  =  8'b00111000;     //97pi/512
  assign sin2[98]  =  8'b11100010;     //98pi/512
  assign cos2[98]  =  8'b00111000;     //98pi/512
  assign sin2[99]  =  8'b11100010;     //99pi/512
  assign cos2[99]  =  8'b00111000;     //99pi/512
  assign sin2[100]  =  8'b11100010;     //100pi/512
  assign cos2[100]  =  8'b00111000;     //100pi/512
  assign sin2[101]  =  8'b11100010;     //101pi/512
  assign cos2[101]  =  8'b00111000;     //101pi/512
  assign sin2[102]  =  8'b11100001;     //102pi/512
  assign cos2[102]  =  8'b00111000;     //102pi/512
  assign sin2[103]  =  8'b11100001;     //103pi/512
  assign cos2[103]  =  8'b00110111;     //103pi/512
  assign sin2[104]  =  8'b11100001;     //104pi/512
  assign cos2[104]  =  8'b00110111;     //104pi/512
  assign sin2[105]  =  8'b11100000;     //105pi/512
  assign cos2[105]  =  8'b00110111;     //105pi/512
  assign sin2[106]  =  8'b11100000;     //106pi/512
  assign cos2[106]  =  8'b00110111;     //106pi/512
  assign sin2[107]  =  8'b11100000;     //107pi/512
  assign cos2[107]  =  8'b00110111;     //107pi/512
  assign sin2[108]  =  8'b11100000;     //108pi/512
  assign cos2[108]  =  8'b00110111;     //108pi/512
  assign sin2[109]  =  8'b11011111;     //109pi/512
  assign cos2[109]  =  8'b00110111;     //109pi/512
  assign sin2[110]  =  8'b11011111;     //110pi/512
  assign cos2[110]  =  8'b00110110;     //110pi/512
  assign sin2[111]  =  8'b11011111;     //111pi/512
  assign cos2[111]  =  8'b00110110;     //111pi/512
  assign sin2[112]  =  8'b11011111;     //112pi/512
  assign cos2[112]  =  8'b00110110;     //112pi/512
  assign sin2[113]  =  8'b11011110;     //113pi/512
  assign cos2[113]  =  8'b00110110;     //113pi/512
  assign sin2[114]  =  8'b11011110;     //114pi/512
  assign cos2[114]  =  8'b00110110;     //114pi/512
  assign sin2[115]  =  8'b11011110;     //115pi/512
  assign cos2[115]  =  8'b00110110;     //115pi/512
  assign sin2[116]  =  8'b11011101;     //116pi/512
  assign cos2[116]  =  8'b00110101;     //116pi/512
  assign sin2[117]  =  8'b11011101;     //117pi/512
  assign cos2[117]  =  8'b00110101;     //117pi/512
  assign sin2[118]  =  8'b11011101;     //118pi/512
  assign cos2[118]  =  8'b00110101;     //118pi/512
  assign sin2[119]  =  8'b11011101;     //119pi/512
  assign cos2[119]  =  8'b00110101;     //119pi/512
  assign sin2[120]  =  8'b11011100;     //120pi/512
  assign cos2[120]  =  8'b00110101;     //120pi/512
  assign sin2[121]  =  8'b11011100;     //121pi/512
  assign cos2[121]  =  8'b00110101;     //121pi/512
  assign sin2[122]  =  8'b11011100;     //122pi/512
  assign cos2[122]  =  8'b00110100;     //122pi/512
  assign sin2[123]  =  8'b11011100;     //123pi/512
  assign cos2[123]  =  8'b00110100;     //123pi/512
  assign sin2[124]  =  8'b11011011;     //124pi/512
  assign cos2[124]  =  8'b00110100;     //124pi/512
  assign sin2[125]  =  8'b11011011;     //125pi/512
  assign cos2[125]  =  8'b00110100;     //125pi/512
  assign sin2[126]  =  8'b11011011;     //126pi/512
  assign cos2[126]  =  8'b00110100;     //126pi/512
  assign sin2[127]  =  8'b11011011;     //127pi/512
  assign cos2[127]  =  8'b00110011;     //127pi/512
  assign sin2[128]  =  8'b11011010;     //128pi/512
  assign cos2[128]  =  8'b00110011;     //128pi/512
  assign sin2[129]  =  8'b11011010;     //129pi/512
  assign cos2[129]  =  8'b00110011;     //129pi/512
  assign sin2[130]  =  8'b11011010;     //130pi/512
  assign cos2[130]  =  8'b00110011;     //130pi/512
  assign sin2[131]  =  8'b11011010;     //131pi/512
  assign cos2[131]  =  8'b00110011;     //131pi/512
  assign sin2[132]  =  8'b11011001;     //132pi/512
  assign cos2[132]  =  8'b00110011;     //132pi/512
  assign sin2[133]  =  8'b11011001;     //133pi/512
  assign cos2[133]  =  8'b00110010;     //133pi/512
  assign sin2[134]  =  8'b11011001;     //134pi/512
  assign cos2[134]  =  8'b00110010;     //134pi/512
  assign sin2[135]  =  8'b11011001;     //135pi/512
  assign cos2[135]  =  8'b00110010;     //135pi/512
  assign sin2[136]  =  8'b11011000;     //136pi/512
  assign cos2[136]  =  8'b00110010;     //136pi/512
  assign sin2[137]  =  8'b11011000;     //137pi/512
  assign cos2[137]  =  8'b00110010;     //137pi/512
  assign sin2[138]  =  8'b11011000;     //138pi/512
  assign cos2[138]  =  8'b00110001;     //138pi/512
  assign sin2[139]  =  8'b11011000;     //139pi/512
  assign cos2[139]  =  8'b00110001;     //139pi/512
  assign sin2[140]  =  8'b11010111;     //140pi/512
  assign cos2[140]  =  8'b00110001;     //140pi/512
  assign sin2[141]  =  8'b11010111;     //141pi/512
  assign cos2[141]  =  8'b00110001;     //141pi/512
  assign sin2[142]  =  8'b11010111;     //142pi/512
  assign cos2[142]  =  8'b00110001;     //142pi/512
  assign sin2[143]  =  8'b11010111;     //143pi/512
  assign cos2[143]  =  8'b00110000;     //143pi/512
  assign sin2[144]  =  8'b11010110;     //144pi/512
  assign cos2[144]  =  8'b00110000;     //144pi/512
  assign sin2[145]  =  8'b11010110;     //145pi/512
  assign cos2[145]  =  8'b00110000;     //145pi/512
  assign sin2[146]  =  8'b11010110;     //146pi/512
  assign cos2[146]  =  8'b00110000;     //146pi/512
  assign sin2[147]  =  8'b11010110;     //147pi/512
  assign cos2[147]  =  8'b00110000;     //147pi/512
  assign sin2[148]  =  8'b11010101;     //148pi/512
  assign cos2[148]  =  8'b00101111;     //148pi/512
  assign sin2[149]  =  8'b11010101;     //149pi/512
  assign cos2[149]  =  8'b00101111;     //149pi/512
  assign sin2[150]  =  8'b11010101;     //150pi/512
  assign cos2[150]  =  8'b00101111;     //150pi/512
  assign sin2[151]  =  8'b11010101;     //151pi/512
  assign cos2[151]  =  8'b00101111;     //151pi/512
  assign sin2[152]  =  8'b11010101;     //152pi/512
  assign cos2[152]  =  8'b00101110;     //152pi/512
  assign sin2[153]  =  8'b11010100;     //153pi/512
  assign cos2[153]  =  8'b00101110;     //153pi/512
  assign sin2[154]  =  8'b11010100;     //154pi/512
  assign cos2[154]  =  8'b00101110;     //154pi/512
  assign sin2[155]  =  8'b11010100;     //155pi/512
  assign cos2[155]  =  8'b00101110;     //155pi/512
  assign sin2[156]  =  8'b11010100;     //156pi/512
  assign cos2[156]  =  8'b00101110;     //156pi/512
  assign sin2[157]  =  8'b11010011;     //157pi/512
  assign cos2[157]  =  8'b00101101;     //157pi/512
  assign sin2[158]  =  8'b11010011;     //158pi/512
  assign cos2[158]  =  8'b00101101;     //158pi/512
  assign sin2[159]  =  8'b11010011;     //159pi/512
  assign cos2[159]  =  8'b00101101;     //159pi/512
  assign sin2[160]  =  8'b11010011;     //160pi/512
  assign cos2[160]  =  8'b00101101;     //160pi/512
  assign sin2[161]  =  8'b11010011;     //161pi/512
  assign cos2[161]  =  8'b00101101;     //161pi/512
  assign sin2[162]  =  8'b11010010;     //162pi/512
  assign cos2[162]  =  8'b00101100;     //162pi/512
  assign sin2[163]  =  8'b11010010;     //163pi/512
  assign cos2[163]  =  8'b00101100;     //163pi/512
  assign sin2[164]  =  8'b11010010;     //164pi/512
  assign cos2[164]  =  8'b00101100;     //164pi/512
  assign sin2[165]  =  8'b11010010;     //165pi/512
  assign cos2[165]  =  8'b00101100;     //165pi/512
  assign sin2[166]  =  8'b11010001;     //166pi/512
  assign cos2[166]  =  8'b00101011;     //166pi/512
  assign sin2[167]  =  8'b11010001;     //167pi/512
  assign cos2[167]  =  8'b00101011;     //167pi/512
  assign sin2[168]  =  8'b11010001;     //168pi/512
  assign cos2[168]  =  8'b00101011;     //168pi/512
  assign sin2[169]  =  8'b11010001;     //169pi/512
  assign cos2[169]  =  8'b00101011;     //169pi/512
  assign sin2[170]  =  8'b11010001;     //170pi/512
  assign cos2[170]  =  8'b00101010;     //170pi/512
  assign sin2[171]  =  8'b11010000;     //171pi/512
  assign cos2[171]  =  8'b00101010;     //171pi/512
  assign sin2[172]  =  8'b11010000;     //172pi/512
  assign cos2[172]  =  8'b00101010;     //172pi/512
  assign sin2[173]  =  8'b11010000;     //173pi/512
  assign cos2[173]  =  8'b00101010;     //173pi/512
  assign sin2[174]  =  8'b11010000;     //174pi/512
  assign cos2[174]  =  8'b00101010;     //174pi/512
  assign sin2[175]  =  8'b11010000;     //175pi/512
  assign cos2[175]  =  8'b00101001;     //175pi/512
  assign sin2[176]  =  8'b11001111;     //176pi/512
  assign cos2[176]  =  8'b00101001;     //176pi/512
  assign sin2[177]  =  8'b11001111;     //177pi/512
  assign cos2[177]  =  8'b00101001;     //177pi/512
  assign sin2[178]  =  8'b11001111;     //178pi/512
  assign cos2[178]  =  8'b00101001;     //178pi/512
  assign sin2[179]  =  8'b11001111;     //179pi/512
  assign cos2[179]  =  8'b00101000;     //179pi/512
  assign sin2[180]  =  8'b11001111;     //180pi/512
  assign cos2[180]  =  8'b00101000;     //180pi/512
  assign sin2[181]  =  8'b11001110;     //181pi/512
  assign cos2[181]  =  8'b00101000;     //181pi/512
  assign sin2[182]  =  8'b11001110;     //182pi/512
  assign cos2[182]  =  8'b00101000;     //182pi/512
  assign sin2[183]  =  8'b11001110;     //183pi/512
  assign cos2[183]  =  8'b00100111;     //183pi/512
  assign sin2[184]  =  8'b11001110;     //184pi/512
  assign cos2[184]  =  8'b00100111;     //184pi/512
  assign sin2[185]  =  8'b11001110;     //185pi/512
  assign cos2[185]  =  8'b00100111;     //185pi/512
  assign sin2[186]  =  8'b11001101;     //186pi/512
  assign cos2[186]  =  8'b00100111;     //186pi/512
  assign sin2[187]  =  8'b11001101;     //187pi/512
  assign cos2[187]  =  8'b00100110;     //187pi/512
  assign sin2[188]  =  8'b11001101;     //188pi/512
  assign cos2[188]  =  8'b00100110;     //188pi/512
  assign sin2[189]  =  8'b11001101;     //189pi/512
  assign cos2[189]  =  8'b00100110;     //189pi/512
  assign sin2[190]  =  8'b11001101;     //190pi/512
  assign cos2[190]  =  8'b00100110;     //190pi/512
  assign sin2[191]  =  8'b11001100;     //191pi/512
  assign cos2[191]  =  8'b00100101;     //191pi/512
  assign sin2[192]  =  8'b11001100;     //192pi/512
  assign cos2[192]  =  8'b00100101;     //192pi/512
  assign sin2[193]  =  8'b11001100;     //193pi/512
  assign cos2[193]  =  8'b00100101;     //193pi/512
  assign sin2[194]  =  8'b11001100;     //194pi/512
  assign cos2[194]  =  8'b00100101;     //194pi/512
  assign sin2[195]  =  8'b11001100;     //195pi/512
  assign cos2[195]  =  8'b00100100;     //195pi/512
  assign sin2[196]  =  8'b11001011;     //196pi/512
  assign cos2[196]  =  8'b00100100;     //196pi/512
  assign sin2[197]  =  8'b11001011;     //197pi/512
  assign cos2[197]  =  8'b00100100;     //197pi/512
  assign sin2[198]  =  8'b11001011;     //198pi/512
  assign cos2[198]  =  8'b00100100;     //198pi/512
  assign sin2[199]  =  8'b11001011;     //199pi/512
  assign cos2[199]  =  8'b00100011;     //199pi/512
  assign sin2[200]  =  8'b11001011;     //200pi/512
  assign cos2[200]  =  8'b00100011;     //200pi/512
  assign sin2[201]  =  8'b11001011;     //201pi/512
  assign cos2[201]  =  8'b00100011;     //201pi/512
  assign sin2[202]  =  8'b11001010;     //202pi/512
  assign cos2[202]  =  8'b00100011;     //202pi/512
  assign sin2[203]  =  8'b11001010;     //203pi/512
  assign cos2[203]  =  8'b00100010;     //203pi/512
  assign sin2[204]  =  8'b11001010;     //204pi/512
  assign cos2[204]  =  8'b00100010;     //204pi/512
  assign sin2[205]  =  8'b11001010;     //205pi/512
  assign cos2[205]  =  8'b00100010;     //205pi/512
  assign sin2[206]  =  8'b11001010;     //206pi/512
  assign cos2[206]  =  8'b00100001;     //206pi/512
  assign sin2[207]  =  8'b11001010;     //207pi/512
  assign cos2[207]  =  8'b00100001;     //207pi/512
  assign sin2[208]  =  8'b11001001;     //208pi/512
  assign cos2[208]  =  8'b00100001;     //208pi/512
  assign sin2[209]  =  8'b11001001;     //209pi/512
  assign cos2[209]  =  8'b00100001;     //209pi/512
  assign sin2[210]  =  8'b11001001;     //210pi/512
  assign cos2[210]  =  8'b00100000;     //210pi/512
  assign sin2[211]  =  8'b11001001;     //211pi/512
  assign cos2[211]  =  8'b00100000;     //211pi/512
  assign sin2[212]  =  8'b11001001;     //212pi/512
  assign cos2[212]  =  8'b00100000;     //212pi/512
  assign sin2[213]  =  8'b11001001;     //213pi/512
  assign cos2[213]  =  8'b00100000;     //213pi/512
  assign sin2[214]  =  8'b11001000;     //214pi/512
  assign cos2[214]  =  8'b00011111;     //214pi/512
  assign sin2[215]  =  8'b11001000;     //215pi/512
  assign cos2[215]  =  8'b00011111;     //215pi/512
  assign sin2[216]  =  8'b11001000;     //216pi/512
  assign cos2[216]  =  8'b00011111;     //216pi/512
  assign sin2[217]  =  8'b11001000;     //217pi/512
  assign cos2[217]  =  8'b00011110;     //217pi/512
  assign sin2[218]  =  8'b11001000;     //218pi/512
  assign cos2[218]  =  8'b00011110;     //218pi/512
  assign sin2[219]  =  8'b11001000;     //219pi/512
  assign cos2[219]  =  8'b00011110;     //219pi/512
  assign sin2[220]  =  8'b11001000;     //220pi/512
  assign cos2[220]  =  8'b00011110;     //220pi/512
  assign sin2[221]  =  8'b11000111;     //221pi/512
  assign cos2[221]  =  8'b00011101;     //221pi/512
  assign sin2[222]  =  8'b11000111;     //222pi/512
  assign cos2[222]  =  8'b00011101;     //222pi/512
  assign sin2[223]  =  8'b11000111;     //223pi/512
  assign cos2[223]  =  8'b00011101;     //223pi/512
  assign sin2[224]  =  8'b11000111;     //224pi/512
  assign cos2[224]  =  8'b00011101;     //224pi/512
  assign sin2[225]  =  8'b11000111;     //225pi/512
  assign cos2[225]  =  8'b00011100;     //225pi/512
  assign sin2[226]  =  8'b11000111;     //226pi/512
  assign cos2[226]  =  8'b00011100;     //226pi/512
  assign sin2[227]  =  8'b11000111;     //227pi/512
  assign cos2[227]  =  8'b00011100;     //227pi/512
  assign sin2[228]  =  8'b11000110;     //228pi/512
  assign cos2[228]  =  8'b00011011;     //228pi/512
  assign sin2[229]  =  8'b11000110;     //229pi/512
  assign cos2[229]  =  8'b00011011;     //229pi/512
  assign sin2[230]  =  8'b11000110;     //230pi/512
  assign cos2[230]  =  8'b00011011;     //230pi/512
  assign sin2[231]  =  8'b11000110;     //231pi/512
  assign cos2[231]  =  8'b00011011;     //231pi/512
  assign sin2[232]  =  8'b11000110;     //232pi/512
  assign cos2[232]  =  8'b00011010;     //232pi/512
  assign sin2[233]  =  8'b11000110;     //233pi/512
  assign cos2[233]  =  8'b00011010;     //233pi/512
  assign sin2[234]  =  8'b11000110;     //234pi/512
  assign cos2[234]  =  8'b00011010;     //234pi/512
  assign sin2[235]  =  8'b11000101;     //235pi/512
  assign cos2[235]  =  8'b00011001;     //235pi/512
  assign sin2[236]  =  8'b11000101;     //236pi/512
  assign cos2[236]  =  8'b00011001;     //236pi/512
  assign sin2[237]  =  8'b11000101;     //237pi/512
  assign cos2[237]  =  8'b00011001;     //237pi/512
  assign sin2[238]  =  8'b11000101;     //238pi/512
  assign cos2[238]  =  8'b00011001;     //238pi/512
  assign sin2[239]  =  8'b11000101;     //239pi/512
  assign cos2[239]  =  8'b00011000;     //239pi/512
  assign sin2[240]  =  8'b11000101;     //240pi/512
  assign cos2[240]  =  8'b00011000;     //240pi/512
  assign sin2[241]  =  8'b11000101;     //241pi/512
  assign cos2[241]  =  8'b00011000;     //241pi/512
  assign sin2[242]  =  8'b11000101;     //242pi/512
  assign cos2[242]  =  8'b00010111;     //242pi/512
  assign sin2[243]  =  8'b11000101;     //243pi/512
  assign cos2[243]  =  8'b00010111;     //243pi/512
  assign sin2[244]  =  8'b11000100;     //244pi/512
  assign cos2[244]  =  8'b00010111;     //244pi/512
  assign sin2[245]  =  8'b11000100;     //245pi/512
  assign cos2[245]  =  8'b00010111;     //245pi/512
  assign sin2[246]  =  8'b11000100;     //246pi/512
  assign cos2[246]  =  8'b00010110;     //246pi/512
  assign sin2[247]  =  8'b11000100;     //247pi/512
  assign cos2[247]  =  8'b00010110;     //247pi/512
  assign sin2[248]  =  8'b11000100;     //248pi/512
  assign cos2[248]  =  8'b00010110;     //248pi/512
  assign sin2[249]  =  8'b11000100;     //249pi/512
  assign cos2[249]  =  8'b00010101;     //249pi/512
  assign sin2[250]  =  8'b11000100;     //250pi/512
  assign cos2[250]  =  8'b00010101;     //250pi/512
  assign sin2[251]  =  8'b11000100;     //251pi/512
  assign cos2[251]  =  8'b00010101;     //251pi/512
  assign sin2[252]  =  8'b11000100;     //252pi/512
  assign cos2[252]  =  8'b00010100;     //252pi/512
  assign sin2[253]  =  8'b11000011;     //253pi/512
  assign cos2[253]  =  8'b00010100;     //253pi/512
  assign sin2[254]  =  8'b11000011;     //254pi/512
  assign cos2[254]  =  8'b00010100;     //254pi/512
  assign sin2[255]  =  8'b11000011;     //255pi/512
  assign cos2[255]  =  8'b00010100;     //255pi/512
  assign sin2[256]  =  8'b11000011;     //256pi/512
  assign cos2[256]  =  8'b00010011;     //256pi/512
  assign sin2[257]  =  8'b11000011;     //257pi/512
  assign cos2[257]  =  8'b00010011;     //257pi/512
  assign sin2[258]  =  8'b11000011;     //258pi/512
  assign cos2[258]  =  8'b00010011;     //258pi/512
  assign sin2[259]  =  8'b11000011;     //259pi/512
  assign cos2[259]  =  8'b00010010;     //259pi/512
  assign sin2[260]  =  8'b11000011;     //260pi/512
  assign cos2[260]  =  8'b00010010;     //260pi/512
  assign sin2[261]  =  8'b11000011;     //261pi/512
  assign cos2[261]  =  8'b00010010;     //261pi/512
  assign sin2[262]  =  8'b11000011;     //262pi/512
  assign cos2[262]  =  8'b00010001;     //262pi/512
  assign sin2[263]  =  8'b11000010;     //263pi/512
  assign cos2[263]  =  8'b00010001;     //263pi/512
  assign sin2[264]  =  8'b11000010;     //264pi/512
  assign cos2[264]  =  8'b00010001;     //264pi/512
  assign sin2[265]  =  8'b11000010;     //265pi/512
  assign cos2[265]  =  8'b00010001;     //265pi/512
  assign sin2[266]  =  8'b11000010;     //266pi/512
  assign cos2[266]  =  8'b00010000;     //266pi/512
  assign sin2[267]  =  8'b11000010;     //267pi/512
  assign cos2[267]  =  8'b00010000;     //267pi/512
  assign sin2[268]  =  8'b11000010;     //268pi/512
  assign cos2[268]  =  8'b00010000;     //268pi/512
  assign sin2[269]  =  8'b11000010;     //269pi/512
  assign cos2[269]  =  8'b00001111;     //269pi/512
  assign sin2[270]  =  8'b11000010;     //270pi/512
  assign cos2[270]  =  8'b00001111;     //270pi/512
  assign sin2[271]  =  8'b11000010;     //271pi/512
  assign cos2[271]  =  8'b00001111;     //271pi/512
  assign sin2[272]  =  8'b11000010;     //272pi/512
  assign cos2[272]  =  8'b00001110;     //272pi/512
  assign sin2[273]  =  8'b11000010;     //273pi/512
  assign cos2[273]  =  8'b00001110;     //273pi/512
  assign sin2[274]  =  8'b11000010;     //274pi/512
  assign cos2[274]  =  8'b00001110;     //274pi/512
  assign sin2[275]  =  8'b11000010;     //275pi/512
  assign cos2[275]  =  8'b00001110;     //275pi/512
  assign sin2[276]  =  8'b11000001;     //276pi/512
  assign cos2[276]  =  8'b00001101;     //276pi/512
  assign sin2[277]  =  8'b11000001;     //277pi/512
  assign cos2[277]  =  8'b00001101;     //277pi/512
  assign sin2[278]  =  8'b11000001;     //278pi/512
  assign cos2[278]  =  8'b00001101;     //278pi/512
  assign sin2[279]  =  8'b11000001;     //279pi/512
  assign cos2[279]  =  8'b00001100;     //279pi/512
  assign sin2[280]  =  8'b11000001;     //280pi/512
  assign cos2[280]  =  8'b00001100;     //280pi/512
  assign sin2[281]  =  8'b11000001;     //281pi/512
  assign cos2[281]  =  8'b00001100;     //281pi/512
  assign sin2[282]  =  8'b11000001;     //282pi/512
  assign cos2[282]  =  8'b00001011;     //282pi/512
  assign sin2[283]  =  8'b11000001;     //283pi/512
  assign cos2[283]  =  8'b00001011;     //283pi/512
  assign sin2[284]  =  8'b11000001;     //284pi/512
  assign cos2[284]  =  8'b00001011;     //284pi/512
  assign sin2[285]  =  8'b11000001;     //285pi/512
  assign cos2[285]  =  8'b00001010;     //285pi/512
  assign sin2[286]  =  8'b11000001;     //286pi/512
  assign cos2[286]  =  8'b00001010;     //286pi/512
  assign sin2[287]  =  8'b11000001;     //287pi/512
  assign cos2[287]  =  8'b00001010;     //287pi/512
  assign sin2[288]  =  8'b11000001;     //288pi/512
  assign cos2[288]  =  8'b00001010;     //288pi/512
  assign sin2[289]  =  8'b11000001;     //289pi/512
  assign cos2[289]  =  8'b00001001;     //289pi/512
  assign sin2[290]  =  8'b11000001;     //290pi/512
  assign cos2[290]  =  8'b00001001;     //290pi/512
  assign sin2[291]  =  8'b11000001;     //291pi/512
  assign cos2[291]  =  8'b00001001;     //291pi/512
  assign sin2[292]  =  8'b11000001;     //292pi/512
  assign cos2[292]  =  8'b00001000;     //292pi/512
  assign sin2[293]  =  8'b11000001;     //293pi/512
  assign cos2[293]  =  8'b00001000;     //293pi/512
  assign sin2[294]  =  8'b11000001;     //294pi/512
  assign cos2[294]  =  8'b00001000;     //294pi/512
  assign sin2[295]  =  8'b11000000;     //295pi/512
  assign cos2[295]  =  8'b00000111;     //295pi/512
  assign sin2[296]  =  8'b11000000;     //296pi/512
  assign cos2[296]  =  8'b00000111;     //296pi/512
  assign sin2[297]  =  8'b11000000;     //297pi/512
  assign cos2[297]  =  8'b00000111;     //297pi/512
  assign sin2[298]  =  8'b11000000;     //298pi/512
  assign cos2[298]  =  8'b00000110;     //298pi/512
  assign sin2[299]  =  8'b11000000;     //299pi/512
  assign cos2[299]  =  8'b00000110;     //299pi/512
  assign sin2[300]  =  8'b11000000;     //300pi/512
  assign cos2[300]  =  8'b00000110;     //300pi/512
  assign sin2[301]  =  8'b11000000;     //301pi/512
  assign cos2[301]  =  8'b00000101;     //301pi/512
  assign sin2[302]  =  8'b11000000;     //302pi/512
  assign cos2[302]  =  8'b00000101;     //302pi/512
  assign sin2[303]  =  8'b11000000;     //303pi/512
  assign cos2[303]  =  8'b00000101;     //303pi/512
  assign sin2[304]  =  8'b11000000;     //304pi/512
  assign cos2[304]  =  8'b00000101;     //304pi/512
  assign sin2[305]  =  8'b11000000;     //305pi/512
  assign cos2[305]  =  8'b00000100;     //305pi/512
  assign sin2[306]  =  8'b11000000;     //306pi/512
  assign cos2[306]  =  8'b00000100;     //306pi/512
  assign sin2[307]  =  8'b11000000;     //307pi/512
  assign cos2[307]  =  8'b00000100;     //307pi/512
  assign sin2[308]  =  8'b11000000;     //308pi/512
  assign cos2[308]  =  8'b00000011;     //308pi/512
  assign sin2[309]  =  8'b11000000;     //309pi/512
  assign cos2[309]  =  8'b00000011;     //309pi/512
  assign sin2[310]  =  8'b11000000;     //310pi/512
  assign cos2[310]  =  8'b00000011;     //310pi/512
  assign sin2[311]  =  8'b11000000;     //311pi/512
  assign cos2[311]  =  8'b00000010;     //311pi/512
  assign sin2[312]  =  8'b11000000;     //312pi/512
  assign cos2[312]  =  8'b00000010;     //312pi/512
  assign sin2[313]  =  8'b11000000;     //313pi/512
  assign cos2[313]  =  8'b00000010;     //313pi/512
  assign sin2[314]  =  8'b11000000;     //314pi/512
  assign cos2[314]  =  8'b00000001;     //314pi/512
  assign sin2[315]  =  8'b11000000;     //315pi/512
  assign cos2[315]  =  8'b00000001;     //315pi/512
  assign sin2[316]  =  8'b11000000;     //316pi/512
  assign cos2[316]  =  8'b00000001;     //316pi/512
  assign sin2[317]  =  8'b11000000;     //317pi/512
  assign cos2[317]  =  8'b00000000;     //317pi/512
  assign sin2[318]  =  8'b11000000;     //318pi/512
  assign cos2[318]  =  8'b00000000;     //318pi/512
  assign sin2[319]  =  8'b11000000;     //319pi/512
  assign cos2[319]  =  8'b00000000;     //319pi/512
  assign sin2[320]  =  8'b11000000;     //320pi/512
  assign cos2[320]  =  8'b00000000;     //320pi/512
  assign sin2[321]  =  8'b11000000;     //321pi/512
  assign cos2[321]  =  8'b00000000;     //321pi/512
  assign sin2[322]  =  8'b11000000;     //322pi/512
  assign cos2[322]  =  8'b11111111;     //322pi/512
  assign sin2[323]  =  8'b11000000;     //323pi/512
  assign cos2[323]  =  8'b11111111;     //323pi/512
  assign sin2[324]  =  8'b11000000;     //324pi/512
  assign cos2[324]  =  8'b11111111;     //324pi/512
  assign sin2[325]  =  8'b11000000;     //325pi/512
  assign cos2[325]  =  8'b11111110;     //325pi/512
  assign sin2[326]  =  8'b11000000;     //326pi/512
  assign cos2[326]  =  8'b11111110;     //326pi/512
  assign sin2[327]  =  8'b11000000;     //327pi/512
  assign cos2[327]  =  8'b11111110;     //327pi/512
  assign sin2[328]  =  8'b11000000;     //328pi/512
  assign cos2[328]  =  8'b11111101;     //328pi/512
  assign sin2[329]  =  8'b11000000;     //329pi/512
  assign cos2[329]  =  8'b11111101;     //329pi/512
  assign sin2[330]  =  8'b11000000;     //330pi/512
  assign cos2[330]  =  8'b11111101;     //330pi/512
  assign sin2[331]  =  8'b11000000;     //331pi/512
  assign cos2[331]  =  8'b11111101;     //331pi/512
  assign sin2[332]  =  8'b11000000;     //332pi/512
  assign cos2[332]  =  8'b11111100;     //332pi/512
  assign sin2[333]  =  8'b11000000;     //333pi/512
  assign cos2[333]  =  8'b11111100;     //333pi/512
  assign sin2[334]  =  8'b11000000;     //334pi/512
  assign cos2[334]  =  8'b11111100;     //334pi/512
  assign sin2[335]  =  8'b11000000;     //335pi/512
  assign cos2[335]  =  8'b11111011;     //335pi/512
  assign sin2[336]  =  8'b11000000;     //336pi/512
  assign cos2[336]  =  8'b11111011;     //336pi/512
  assign sin2[337]  =  8'b11000000;     //337pi/512
  assign cos2[337]  =  8'b11111011;     //337pi/512
  assign sin2[338]  =  8'b11000000;     //338pi/512
  assign cos2[338]  =  8'b11111010;     //338pi/512
  assign sin2[339]  =  8'b11000000;     //339pi/512
  assign cos2[339]  =  8'b11111010;     //339pi/512
  assign sin2[340]  =  8'b11000000;     //340pi/512
  assign cos2[340]  =  8'b11111010;     //340pi/512
  assign sin2[341]  =  8'b11000000;     //341pi/512
  assign cos2[341]  =  8'b11111001;     //341pi/512
  assign sin2[342]  =  8'b11000000;     //342pi/512
  assign cos2[342]  =  8'b11111001;     //342pi/512
  assign sin2[343]  =  8'b11000000;     //343pi/512
  assign cos2[343]  =  8'b11111001;     //343pi/512
  assign sin2[344]  =  8'b11000000;     //344pi/512
  assign cos2[344]  =  8'b11111000;     //344pi/512
  assign sin2[345]  =  8'b11000000;     //345pi/512
  assign cos2[345]  =  8'b11111000;     //345pi/512
  assign sin2[346]  =  8'b11000001;     //346pi/512
  assign cos2[346]  =  8'b11111000;     //346pi/512
  assign sin2[347]  =  8'b11000001;     //347pi/512
  assign cos2[347]  =  8'b11111000;     //347pi/512
  assign sin2[348]  =  8'b11000001;     //348pi/512
  assign cos2[348]  =  8'b11110111;     //348pi/512
  assign sin2[349]  =  8'b11000001;     //349pi/512
  assign cos2[349]  =  8'b11110111;     //349pi/512
  assign sin2[350]  =  8'b11000001;     //350pi/512
  assign cos2[350]  =  8'b11110111;     //350pi/512
  assign sin2[351]  =  8'b11000001;     //351pi/512
  assign cos2[351]  =  8'b11110110;     //351pi/512
  assign sin2[352]  =  8'b11000001;     //352pi/512
  assign cos2[352]  =  8'b11110110;     //352pi/512
  assign sin2[353]  =  8'b11000001;     //353pi/512
  assign cos2[353]  =  8'b11110110;     //353pi/512
  assign sin2[354]  =  8'b11000001;     //354pi/512
  assign cos2[354]  =  8'b11110101;     //354pi/512
  assign sin2[355]  =  8'b11000001;     //355pi/512
  assign cos2[355]  =  8'b11110101;     //355pi/512
  assign sin2[356]  =  8'b11000001;     //356pi/512
  assign cos2[356]  =  8'b11110101;     //356pi/512
  assign sin2[357]  =  8'b11000001;     //357pi/512
  assign cos2[357]  =  8'b11110100;     //357pi/512
  assign sin2[358]  =  8'b11000001;     //358pi/512
  assign cos2[358]  =  8'b11110100;     //358pi/512
  assign sin2[359]  =  8'b11000001;     //359pi/512
  assign cos2[359]  =  8'b11110100;     //359pi/512
  assign sin2[360]  =  8'b11000001;     //360pi/512
  assign cos2[360]  =  8'b11110100;     //360pi/512
  assign sin2[361]  =  8'b11000001;     //361pi/512
  assign cos2[361]  =  8'b11110011;     //361pi/512
  assign sin2[362]  =  8'b11000001;     //362pi/512
  assign cos2[362]  =  8'b11110011;     //362pi/512
  assign sin2[363]  =  8'b11000001;     //363pi/512
  assign cos2[363]  =  8'b11110011;     //363pi/512
  assign sin2[364]  =  8'b11000001;     //364pi/512
  assign cos2[364]  =  8'b11110010;     //364pi/512
  assign sin2[365]  =  8'b11000010;     //365pi/512
  assign cos2[365]  =  8'b11110010;     //365pi/512
  assign sin2[366]  =  8'b11000010;     //366pi/512
  assign cos2[366]  =  8'b11110010;     //366pi/512
  assign sin2[367]  =  8'b11000010;     //367pi/512
  assign cos2[367]  =  8'b11110001;     //367pi/512
  assign sin2[368]  =  8'b11000010;     //368pi/512
  assign cos2[368]  =  8'b11110001;     //368pi/512
  assign sin2[369]  =  8'b11000010;     //369pi/512
  assign cos2[369]  =  8'b11110001;     //369pi/512
  assign sin2[370]  =  8'b11000010;     //370pi/512
  assign cos2[370]  =  8'b11110000;     //370pi/512
  assign sin2[371]  =  8'b11000010;     //371pi/512
  assign cos2[371]  =  8'b11110000;     //371pi/512
  assign sin2[372]  =  8'b11000010;     //372pi/512
  assign cos2[372]  =  8'b11110000;     //372pi/512
  assign sin2[373]  =  8'b11000010;     //373pi/512
  assign cos2[373]  =  8'b11110000;     //373pi/512
  assign sin2[374]  =  8'b11000010;     //374pi/512
  assign cos2[374]  =  8'b11101111;     //374pi/512
  assign sin2[375]  =  8'b11000010;     //375pi/512
  assign cos2[375]  =  8'b11101111;     //375pi/512
  assign sin2[376]  =  8'b11000010;     //376pi/512
  assign cos2[376]  =  8'b11101111;     //376pi/512
  assign sin2[377]  =  8'b11000010;     //377pi/512
  assign cos2[377]  =  8'b11101110;     //377pi/512
  assign sin2[378]  =  8'b11000011;     //378pi/512
  assign cos2[378]  =  8'b11101110;     //378pi/512
  assign sin2[379]  =  8'b11000011;     //379pi/512
  assign cos2[379]  =  8'b11101110;     //379pi/512
  assign sin2[380]  =  8'b11000011;     //380pi/512
  assign cos2[380]  =  8'b11101101;     //380pi/512
  assign sin2[381]  =  8'b11000011;     //381pi/512
  assign cos2[381]  =  8'b11101101;     //381pi/512
  assign sin2[382]  =  8'b11000011;     //382pi/512
  assign cos2[382]  =  8'b11101101;     //382pi/512
  assign sin2[383]  =  8'b11000011;     //383pi/512
  assign cos2[383]  =  8'b11101101;     //383pi/512
  assign sin2[384]  =  8'b11000011;     //384pi/512
  assign cos2[384]  =  8'b11101100;     //384pi/512
  assign sin2[385]  =  8'b11000011;     //385pi/512
  assign cos2[385]  =  8'b11101100;     //385pi/512
  assign sin2[386]  =  8'b11000011;     //386pi/512
  assign cos2[386]  =  8'b11101100;     //386pi/512
  assign sin2[387]  =  8'b11000011;     //387pi/512
  assign cos2[387]  =  8'b11101011;     //387pi/512
  assign sin2[388]  =  8'b11000100;     //388pi/512
  assign cos2[388]  =  8'b11101011;     //388pi/512
  assign sin2[389]  =  8'b11000100;     //389pi/512
  assign cos2[389]  =  8'b11101011;     //389pi/512
  assign sin2[390]  =  8'b11000100;     //390pi/512
  assign cos2[390]  =  8'b11101010;     //390pi/512
  assign sin2[391]  =  8'b11000100;     //391pi/512
  assign cos2[391]  =  8'b11101010;     //391pi/512
  assign sin2[392]  =  8'b11000100;     //392pi/512
  assign cos2[392]  =  8'b11101010;     //392pi/512
  assign sin2[393]  =  8'b11000100;     //393pi/512
  assign cos2[393]  =  8'b11101010;     //393pi/512
  assign sin2[394]  =  8'b11000100;     //394pi/512
  assign cos2[394]  =  8'b11101001;     //394pi/512
  assign sin2[395]  =  8'b11000100;     //395pi/512
  assign cos2[395]  =  8'b11101001;     //395pi/512
  assign sin2[396]  =  8'b11000100;     //396pi/512
  assign cos2[396]  =  8'b11101001;     //396pi/512
  assign sin2[397]  =  8'b11000101;     //397pi/512
  assign cos2[397]  =  8'b11101000;     //397pi/512
  assign sin2[398]  =  8'b11000101;     //398pi/512
  assign cos2[398]  =  8'b11101000;     //398pi/512
  assign sin2[399]  =  8'b11000101;     //399pi/512
  assign cos2[399]  =  8'b11101000;     //399pi/512
  assign sin2[400]  =  8'b11000101;     //400pi/512
  assign cos2[400]  =  8'b11101000;     //400pi/512
  assign sin2[401]  =  8'b11000101;     //401pi/512
  assign cos2[401]  =  8'b11100111;     //401pi/512
  assign sin2[402]  =  8'b11000101;     //402pi/512
  assign cos2[402]  =  8'b11100111;     //402pi/512
  assign sin2[403]  =  8'b11000101;     //403pi/512
  assign cos2[403]  =  8'b11100111;     //403pi/512
  assign sin2[404]  =  8'b11000101;     //404pi/512
  assign cos2[404]  =  8'b11100110;     //404pi/512
  assign sin2[405]  =  8'b11000101;     //405pi/512
  assign cos2[405]  =  8'b11100110;     //405pi/512
  assign sin2[406]  =  8'b11000110;     //406pi/512
  assign cos2[406]  =  8'b11100110;     //406pi/512
  assign sin2[407]  =  8'b11000110;     //407pi/512
  assign cos2[407]  =  8'b11100101;     //407pi/512
  assign sin2[408]  =  8'b11000110;     //408pi/512
  assign cos2[408]  =  8'b11100101;     //408pi/512
  assign sin2[409]  =  8'b11000110;     //409pi/512
  assign cos2[409]  =  8'b11100101;     //409pi/512
  assign sin2[410]  =  8'b11000110;     //410pi/512
  assign cos2[410]  =  8'b11100101;     //410pi/512
  assign sin2[411]  =  8'b11000110;     //411pi/512
  assign cos2[411]  =  8'b11100100;     //411pi/512
  assign sin2[412]  =  8'b11000110;     //412pi/512
  assign cos2[412]  =  8'b11100100;     //412pi/512
  assign sin2[413]  =  8'b11000111;     //413pi/512
  assign cos2[413]  =  8'b11100100;     //413pi/512
  assign sin2[414]  =  8'b11000111;     //414pi/512
  assign cos2[414]  =  8'b11100100;     //414pi/512
  assign sin2[415]  =  8'b11000111;     //415pi/512
  assign cos2[415]  =  8'b11100011;     //415pi/512
  assign sin2[416]  =  8'b11000111;     //416pi/512
  assign cos2[416]  =  8'b11100011;     //416pi/512
  assign sin2[417]  =  8'b11000111;     //417pi/512
  assign cos2[417]  =  8'b11100011;     //417pi/512
  assign sin2[418]  =  8'b11000111;     //418pi/512
  assign cos2[418]  =  8'b11100010;     //418pi/512
  assign sin2[419]  =  8'b11000111;     //419pi/512
  assign cos2[419]  =  8'b11100010;     //419pi/512
  assign sin2[420]  =  8'b11001000;     //420pi/512
  assign cos2[420]  =  8'b11100010;     //420pi/512
  assign sin2[421]  =  8'b11001000;     //421pi/512
  assign cos2[421]  =  8'b11100010;     //421pi/512
  assign sin2[422]  =  8'b11001000;     //422pi/512
  assign cos2[422]  =  8'b11100001;     //422pi/512
  assign sin2[423]  =  8'b11001000;     //423pi/512
  assign cos2[423]  =  8'b11100001;     //423pi/512
  assign sin2[424]  =  8'b11001000;     //424pi/512
  assign cos2[424]  =  8'b11100001;     //424pi/512
  assign sin2[425]  =  8'b11001000;     //425pi/512
  assign cos2[425]  =  8'b11100000;     //425pi/512
  assign sin2[426]  =  8'b11001000;     //426pi/512
  assign cos2[426]  =  8'b11100000;     //426pi/512
  assign sin2[427]  =  8'b11001001;     //427pi/512
  assign cos2[427]  =  8'b11100000;     //427pi/512
  assign sin2[428]  =  8'b11001001;     //428pi/512
  assign cos2[428]  =  8'b11100000;     //428pi/512
  assign sin2[429]  =  8'b11001001;     //429pi/512
  assign cos2[429]  =  8'b11011111;     //429pi/512
  assign sin2[430]  =  8'b11001001;     //430pi/512
  assign cos2[430]  =  8'b11011111;     //430pi/512
  assign sin2[431]  =  8'b11001001;     //431pi/512
  assign cos2[431]  =  8'b11011111;     //431pi/512
  assign sin2[432]  =  8'b11001001;     //432pi/512
  assign cos2[432]  =  8'b11011111;     //432pi/512
  assign sin2[433]  =  8'b11001010;     //433pi/512
  assign cos2[433]  =  8'b11011110;     //433pi/512
  assign sin2[434]  =  8'b11001010;     //434pi/512
  assign cos2[434]  =  8'b11011110;     //434pi/512
  assign sin2[435]  =  8'b11001010;     //435pi/512
  assign cos2[435]  =  8'b11011110;     //435pi/512
  assign sin2[436]  =  8'b11001010;     //436pi/512
  assign cos2[436]  =  8'b11011101;     //436pi/512
  assign sin2[437]  =  8'b11001010;     //437pi/512
  assign cos2[437]  =  8'b11011101;     //437pi/512
  assign sin2[438]  =  8'b11001010;     //438pi/512
  assign cos2[438]  =  8'b11011101;     //438pi/512
  assign sin2[439]  =  8'b11001011;     //439pi/512
  assign cos2[439]  =  8'b11011101;     //439pi/512
  assign sin2[440]  =  8'b11001011;     //440pi/512
  assign cos2[440]  =  8'b11011100;     //440pi/512
  assign sin2[441]  =  8'b11001011;     //441pi/512
  assign cos2[441]  =  8'b11011100;     //441pi/512
  assign sin2[442]  =  8'b11001011;     //442pi/512
  assign cos2[442]  =  8'b11011100;     //442pi/512
  assign sin2[443]  =  8'b11001011;     //443pi/512
  assign cos2[443]  =  8'b11011100;     //443pi/512
  assign sin2[444]  =  8'b11001011;     //444pi/512
  assign cos2[444]  =  8'b11011011;     //444pi/512
  assign sin2[445]  =  8'b11001100;     //445pi/512
  assign cos2[445]  =  8'b11011011;     //445pi/512
  assign sin2[446]  =  8'b11001100;     //446pi/512
  assign cos2[446]  =  8'b11011011;     //446pi/512
  assign sin2[447]  =  8'b11001100;     //447pi/512
  assign cos2[447]  =  8'b11011011;     //447pi/512
  assign sin2[448]  =  8'b11001100;     //448pi/512
  assign cos2[448]  =  8'b11011010;     //448pi/512
  assign sin2[449]  =  8'b11001100;     //449pi/512
  assign cos2[449]  =  8'b11011010;     //449pi/512
  assign sin2[450]  =  8'b11001101;     //450pi/512
  assign cos2[450]  =  8'b11011010;     //450pi/512
  assign sin2[451]  =  8'b11001101;     //451pi/512
  assign cos2[451]  =  8'b11011010;     //451pi/512
  assign sin2[452]  =  8'b11001101;     //452pi/512
  assign cos2[452]  =  8'b11011001;     //452pi/512
  assign sin2[453]  =  8'b11001101;     //453pi/512
  assign cos2[453]  =  8'b11011001;     //453pi/512
  assign sin2[454]  =  8'b11001101;     //454pi/512
  assign cos2[454]  =  8'b11011001;     //454pi/512
  assign sin2[455]  =  8'b11001110;     //455pi/512
  assign cos2[455]  =  8'b11011001;     //455pi/512
  assign sin2[456]  =  8'b11001110;     //456pi/512
  assign cos2[456]  =  8'b11011000;     //456pi/512
  assign sin2[457]  =  8'b11001110;     //457pi/512
  assign cos2[457]  =  8'b11011000;     //457pi/512
  assign sin2[458]  =  8'b11001110;     //458pi/512
  assign cos2[458]  =  8'b11011000;     //458pi/512
  assign sin2[459]  =  8'b11001110;     //459pi/512
  assign cos2[459]  =  8'b11011000;     //459pi/512
  assign sin2[460]  =  8'b11001111;     //460pi/512
  assign cos2[460]  =  8'b11010111;     //460pi/512
  assign sin2[461]  =  8'b11001111;     //461pi/512
  assign cos2[461]  =  8'b11010111;     //461pi/512
  assign sin2[462]  =  8'b11001111;     //462pi/512
  assign cos2[462]  =  8'b11010111;     //462pi/512
  assign sin2[463]  =  8'b11001111;     //463pi/512
  assign cos2[463]  =  8'b11010111;     //463pi/512
  assign sin2[464]  =  8'b11001111;     //464pi/512
  assign cos2[464]  =  8'b11010110;     //464pi/512
  assign sin2[465]  =  8'b11010000;     //465pi/512
  assign cos2[465]  =  8'b11010110;     //465pi/512
  assign sin2[466]  =  8'b11010000;     //466pi/512
  assign cos2[466]  =  8'b11010110;     //466pi/512
  assign sin2[467]  =  8'b11010000;     //467pi/512
  assign cos2[467]  =  8'b11010110;     //467pi/512
  assign sin2[468]  =  8'b11010000;     //468pi/512
  assign cos2[468]  =  8'b11010101;     //468pi/512
  assign sin2[469]  =  8'b11010000;     //469pi/512
  assign cos2[469]  =  8'b11010101;     //469pi/512
  assign sin2[470]  =  8'b11010001;     //470pi/512
  assign cos2[470]  =  8'b11010101;     //470pi/512
  assign sin2[471]  =  8'b11010001;     //471pi/512
  assign cos2[471]  =  8'b11010101;     //471pi/512
  assign sin2[472]  =  8'b11010001;     //472pi/512
  assign cos2[472]  =  8'b11010101;     //472pi/512
  assign sin2[473]  =  8'b11010001;     //473pi/512
  assign cos2[473]  =  8'b11010100;     //473pi/512
  assign sin2[474]  =  8'b11010001;     //474pi/512
  assign cos2[474]  =  8'b11010100;     //474pi/512
  assign sin2[475]  =  8'b11010010;     //475pi/512
  assign cos2[475]  =  8'b11010100;     //475pi/512
  assign sin2[476]  =  8'b11010010;     //476pi/512
  assign cos2[476]  =  8'b11010100;     //476pi/512
  assign sin2[477]  =  8'b11010010;     //477pi/512
  assign cos2[477]  =  8'b11010011;     //477pi/512
  assign sin2[478]  =  8'b11010010;     //478pi/512
  assign cos2[478]  =  8'b11010011;     //478pi/512
  assign sin2[479]  =  8'b11010011;     //479pi/512
  assign cos2[479]  =  8'b11010011;     //479pi/512
  assign sin2[480]  =  8'b11010011;     //480pi/512
  assign cos2[480]  =  8'b11010011;     //480pi/512
  assign sin2[481]  =  8'b11010011;     //481pi/512
  assign cos2[481]  =  8'b11010011;     //481pi/512
  assign sin2[482]  =  8'b11010011;     //482pi/512
  assign cos2[482]  =  8'b11010010;     //482pi/512
  assign sin2[483]  =  8'b11010011;     //483pi/512
  assign cos2[483]  =  8'b11010010;     //483pi/512
  assign sin2[484]  =  8'b11010100;     //484pi/512
  assign cos2[484]  =  8'b11010010;     //484pi/512
  assign sin2[485]  =  8'b11010100;     //485pi/512
  assign cos2[485]  =  8'b11010010;     //485pi/512
  assign sin2[486]  =  8'b11010100;     //486pi/512
  assign cos2[486]  =  8'b11010001;     //486pi/512
  assign sin2[487]  =  8'b11010100;     //487pi/512
  assign cos2[487]  =  8'b11010001;     //487pi/512
  assign sin2[488]  =  8'b11010101;     //488pi/512
  assign cos2[488]  =  8'b11010001;     //488pi/512
  assign sin2[489]  =  8'b11010101;     //489pi/512
  assign cos2[489]  =  8'b11010001;     //489pi/512
  assign sin2[490]  =  8'b11010101;     //490pi/512
  assign cos2[490]  =  8'b11010001;     //490pi/512
  assign sin2[491]  =  8'b11010101;     //491pi/512
  assign cos2[491]  =  8'b11010000;     //491pi/512
  assign sin2[492]  =  8'b11010101;     //492pi/512
  assign cos2[492]  =  8'b11010000;     //492pi/512
  assign sin2[493]  =  8'b11010110;     //493pi/512
  assign cos2[493]  =  8'b11010000;     //493pi/512
  assign sin2[494]  =  8'b11010110;     //494pi/512
  assign cos2[494]  =  8'b11010000;     //494pi/512
  assign sin2[495]  =  8'b11010110;     //495pi/512
  assign cos2[495]  =  8'b11010000;     //495pi/512
  assign sin2[496]  =  8'b11010110;     //496pi/512
  assign cos2[496]  =  8'b11001111;     //496pi/512
  assign sin2[497]  =  8'b11010111;     //497pi/512
  assign cos2[497]  =  8'b11001111;     //497pi/512
  assign sin2[498]  =  8'b11010111;     //498pi/512
  assign cos2[498]  =  8'b11001111;     //498pi/512
  assign sin2[499]  =  8'b11010111;     //499pi/512
  assign cos2[499]  =  8'b11001111;     //499pi/512
  assign sin2[500]  =  8'b11010111;     //500pi/512
  assign cos2[500]  =  8'b11001111;     //500pi/512
  assign sin2[501]  =  8'b11011000;     //501pi/512
  assign cos2[501]  =  8'b11001110;     //501pi/512
  assign sin2[502]  =  8'b11011000;     //502pi/512
  assign cos2[502]  =  8'b11001110;     //502pi/512
  assign sin2[503]  =  8'b11011000;     //503pi/512
  assign cos2[503]  =  8'b11001110;     //503pi/512
  assign sin2[504]  =  8'b11011000;     //504pi/512
  assign cos2[504]  =  8'b11001110;     //504pi/512
  assign sin2[505]  =  8'b11011001;     //505pi/512
  assign cos2[505]  =  8'b11001110;     //505pi/512
  assign sin2[506]  =  8'b11011001;     //506pi/512
  assign cos2[506]  =  8'b11001101;     //506pi/512
  assign sin2[507]  =  8'b11011001;     //507pi/512
  assign cos2[507]  =  8'b11001101;     //507pi/512
  assign sin2[508]  =  8'b11011001;     //508pi/512
  assign cos2[508]  =  8'b11001101;     //508pi/512
  assign sin2[509]  =  8'b11011010;     //509pi/512
  assign cos2[509]  =  8'b11001101;     //509pi/512
  assign sin2[510]  =  8'b11011010;     //510pi/512
  assign cos2[510]  =  8'b11001101;     //510pi/512
  assign sin2[511]  =  8'b11011010;     //511pi/512
  assign cos2[511]  =  8'b11001100;     //511pi/512
 
endmodule