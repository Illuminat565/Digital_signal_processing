module  M_TWIDLE_7_bit #(parameter SIZE =10, word_length_tw = 7) (
    input            clk,
    input            en_rd, 
    input   [10:0]   rd_ptr_angle,
    input            en_modf, 

    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );


reg signed [word_length_tw-1:0]  cos  [511:0];
reg signed [word_length_tw-1:0]  sin  [511:0];

reg signed [word_length_tw-1:0]  m_cos  [511:0];
reg signed [word_length_tw-1:0]  m_sin  [511:0];

reg signed [word_length_tw-1:0]  cos_temp;
reg signed [word_length_tw-1:0]  sin_temp;

reg signed [word_length_tw-1:0]  m_cos_temp;
reg signed [word_length_tw-1:0]  m_sin_temp;


//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & ~ en_modf ) begin
                  cos_temp           <= cos   [rd_ptr_angle];
                  sin_temp           <= sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & en_modf ) begin
                  m_cos_temp           <= m_cos   [rd_ptr_angle];
                  m_sin_temp           <= m_sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(*) begin 
             if (en_modf ) begin
                  cos_data           <= m_cos_temp;
                  sin_data           <= m_sin_temp;
             end else begin
                  cos_data           <= cos_temp;
                  sin_data           <= sin_temp;
             end
        end
//----------------------------------------------------------------------------------------
initial begin

   sin[0]  =  7'b0000000;     //0pi/512
   cos[0]  =  7'b0100000;     //0pi/512
   sin[1]  =  7'b0000000;     //1pi/512
   cos[1]  =  7'b0011111;     //1pi/512
   sin[2]  =  7'b0000000;     //2pi/512
   cos[2]  =  7'b0011111;     //2pi/512
   sin[3]  =  7'b1111111;     //3pi/512
   cos[3]  =  7'b0011111;     //3pi/512
   sin[4]  =  7'b1111111;     //4pi/512
   cos[4]  =  7'b0011111;     //4pi/512
   sin[5]  =  7'b1111111;     //5pi/512
   cos[5]  =  7'b0011111;     //5pi/512
   sin[6]  =  7'b1111111;     //6pi/512
   cos[6]  =  7'b0011111;     //6pi/512
   sin[7]  =  7'b1111111;     //7pi/512
   cos[7]  =  7'b0011111;     //7pi/512
   sin[8]  =  7'b1111110;     //8pi/512
   cos[8]  =  7'b0011111;     //8pi/512
   sin[9]  =  7'b1111110;     //9pi/512
   cos[9]  =  7'b0011111;     //9pi/512
   sin[10]  =  7'b1111110;     //10pi/512
   cos[10]  =  7'b0011111;     //10pi/512
   sin[11]  =  7'b1111110;     //11pi/512
   cos[11]  =  7'b0011111;     //11pi/512
   sin[12]  =  7'b1111110;     //12pi/512
   cos[12]  =  7'b0011111;     //12pi/512
   sin[13]  =  7'b1111101;     //13pi/512
   cos[13]  =  7'b0011111;     //13pi/512
   sin[14]  =  7'b1111101;     //14pi/512
   cos[14]  =  7'b0011111;     //14pi/512
   sin[15]  =  7'b1111101;     //15pi/512
   cos[15]  =  7'b0011111;     //15pi/512
   sin[16]  =  7'b1111101;     //16pi/512
   cos[16]  =  7'b0011111;     //16pi/512
   sin[17]  =  7'b1111101;     //17pi/512
   cos[17]  =  7'b0011111;     //17pi/512
   sin[18]  =  7'b1111100;     //18pi/512
   cos[18]  =  7'b0011111;     //18pi/512
   sin[19]  =  7'b1111100;     //19pi/512
   cos[19]  =  7'b0011111;     //19pi/512
   sin[20]  =  7'b1111100;     //20pi/512
   cos[20]  =  7'b0011111;     //20pi/512
   sin[21]  =  7'b1111100;     //21pi/512
   cos[21]  =  7'b0011111;     //21pi/512
   sin[22]  =  7'b1111100;     //22pi/512
   cos[22]  =  7'b0011111;     //22pi/512
   sin[23]  =  7'b1111011;     //23pi/512
   cos[23]  =  7'b0011111;     //23pi/512
   sin[24]  =  7'b1111011;     //24pi/512
   cos[24]  =  7'b0011111;     //24pi/512
   sin[25]  =  7'b1111011;     //25pi/512
   cos[25]  =  7'b0011111;     //25pi/512
   sin[26]  =  7'b1111011;     //26pi/512
   cos[26]  =  7'b0011111;     //26pi/512
   sin[27]  =  7'b1111011;     //27pi/512
   cos[27]  =  7'b0011111;     //27pi/512
   sin[28]  =  7'b1111011;     //28pi/512
   cos[28]  =  7'b0011111;     //28pi/512
   sin[29]  =  7'b1111010;     //29pi/512
   cos[29]  =  7'b0011111;     //29pi/512
   sin[30]  =  7'b1111010;     //30pi/512
   cos[30]  =  7'b0011111;     //30pi/512
   sin[31]  =  7'b1111010;     //31pi/512
   cos[31]  =  7'b0011111;     //31pi/512
   sin[32]  =  7'b1111010;     //32pi/512
   cos[32]  =  7'b0011111;     //32pi/512
   sin[33]  =  7'b1111010;     //33pi/512
   cos[33]  =  7'b0011111;     //33pi/512
   sin[34]  =  7'b1111001;     //34pi/512
   cos[34]  =  7'b0011111;     //34pi/512
   sin[35]  =  7'b1111001;     //35pi/512
   cos[35]  =  7'b0011111;     //35pi/512
   sin[36]  =  7'b1111001;     //36pi/512
   cos[36]  =  7'b0011111;     //36pi/512
   sin[37]  =  7'b1111001;     //37pi/512
   cos[37]  =  7'b0011111;     //37pi/512
   sin[38]  =  7'b1111001;     //38pi/512
   cos[38]  =  7'b0011111;     //38pi/512
   sin[39]  =  7'b1111000;     //39pi/512
   cos[39]  =  7'b0011111;     //39pi/512
   sin[40]  =  7'b1111000;     //40pi/512
   cos[40]  =  7'b0011111;     //40pi/512
   sin[41]  =  7'b1111000;     //41pi/512
   cos[41]  =  7'b0011110;     //41pi/512
   sin[42]  =  7'b1111000;     //42pi/512
   cos[42]  =  7'b0011110;     //42pi/512
   sin[43]  =  7'b1111000;     //43pi/512
   cos[43]  =  7'b0011110;     //43pi/512
   sin[44]  =  7'b1110111;     //44pi/512
   cos[44]  =  7'b0011110;     //44pi/512
   sin[45]  =  7'b1110111;     //45pi/512
   cos[45]  =  7'b0011110;     //45pi/512
   sin[46]  =  7'b1110111;     //46pi/512
   cos[46]  =  7'b0011110;     //46pi/512
   sin[47]  =  7'b1110111;     //47pi/512
   cos[47]  =  7'b0011110;     //47pi/512
   sin[48]  =  7'b1110111;     //48pi/512
   cos[48]  =  7'b0011110;     //48pi/512
   sin[49]  =  7'b1110111;     //49pi/512
   cos[49]  =  7'b0011110;     //49pi/512
   sin[50]  =  7'b1110110;     //50pi/512
   cos[50]  =  7'b0011110;     //50pi/512
   sin[51]  =  7'b1110110;     //51pi/512
   cos[51]  =  7'b0011110;     //51pi/512
   sin[52]  =  7'b1110110;     //52pi/512
   cos[52]  =  7'b0011110;     //52pi/512
   sin[53]  =  7'b1110110;     //53pi/512
   cos[53]  =  7'b0011110;     //53pi/512
   sin[54]  =  7'b1110110;     //54pi/512
   cos[54]  =  7'b0011110;     //54pi/512
   sin[55]  =  7'b1110101;     //55pi/512
   cos[55]  =  7'b0011110;     //55pi/512
   sin[56]  =  7'b1110101;     //56pi/512
   cos[56]  =  7'b0011110;     //56pi/512
   sin[57]  =  7'b1110101;     //57pi/512
   cos[57]  =  7'b0011110;     //57pi/512
   sin[58]  =  7'b1110101;     //58pi/512
   cos[58]  =  7'b0011101;     //58pi/512
   sin[59]  =  7'b1110101;     //59pi/512
   cos[59]  =  7'b0011101;     //59pi/512
   sin[60]  =  7'b1110100;     //60pi/512
   cos[60]  =  7'b0011101;     //60pi/512
   sin[61]  =  7'b1110100;     //61pi/512
   cos[61]  =  7'b0011101;     //61pi/512
   sin[62]  =  7'b1110100;     //62pi/512
   cos[62]  =  7'b0011101;     //62pi/512
   sin[63]  =  7'b1110100;     //63pi/512
   cos[63]  =  7'b0011101;     //63pi/512
   sin[64]  =  7'b1110100;     //64pi/512
   cos[64]  =  7'b0011101;     //64pi/512
   sin[65]  =  7'b1110100;     //65pi/512
   cos[65]  =  7'b0011101;     //65pi/512
   sin[66]  =  7'b1110011;     //66pi/512
   cos[66]  =  7'b0011101;     //66pi/512
   sin[67]  =  7'b1110011;     //67pi/512
   cos[67]  =  7'b0011101;     //67pi/512
   sin[68]  =  7'b1110011;     //68pi/512
   cos[68]  =  7'b0011101;     //68pi/512
   sin[69]  =  7'b1110011;     //69pi/512
   cos[69]  =  7'b0011101;     //69pi/512
   sin[70]  =  7'b1110011;     //70pi/512
   cos[70]  =  7'b0011101;     //70pi/512
   sin[71]  =  7'b1110010;     //71pi/512
   cos[71]  =  7'b0011101;     //71pi/512
   sin[72]  =  7'b1110010;     //72pi/512
   cos[72]  =  7'b0011100;     //72pi/512
   sin[73]  =  7'b1110010;     //73pi/512
   cos[73]  =  7'b0011100;     //73pi/512
   sin[74]  =  7'b1110010;     //74pi/512
   cos[74]  =  7'b0011100;     //74pi/512
   sin[75]  =  7'b1110010;     //75pi/512
   cos[75]  =  7'b0011100;     //75pi/512
   sin[76]  =  7'b1110010;     //76pi/512
   cos[76]  =  7'b0011100;     //76pi/512
   sin[77]  =  7'b1110001;     //77pi/512
   cos[77]  =  7'b0011100;     //77pi/512
   sin[78]  =  7'b1110001;     //78pi/512
   cos[78]  =  7'b0011100;     //78pi/512
   sin[79]  =  7'b1110001;     //79pi/512
   cos[79]  =  7'b0011100;     //79pi/512
   sin[80]  =  7'b1110001;     //80pi/512
   cos[80]  =  7'b0011100;     //80pi/512
   sin[81]  =  7'b1110001;     //81pi/512
   cos[81]  =  7'b0011100;     //81pi/512
   sin[82]  =  7'b1110001;     //82pi/512
   cos[82]  =  7'b0011100;     //82pi/512
   sin[83]  =  7'b1110000;     //83pi/512
   cos[83]  =  7'b0011011;     //83pi/512
   sin[84]  =  7'b1110000;     //84pi/512
   cos[84]  =  7'b0011011;     //84pi/512
   sin[85]  =  7'b1110000;     //85pi/512
   cos[85]  =  7'b0011011;     //85pi/512
   sin[86]  =  7'b1110000;     //86pi/512
   cos[86]  =  7'b0011011;     //86pi/512
   sin[87]  =  7'b1110000;     //87pi/512
   cos[87]  =  7'b0011011;     //87pi/512
   sin[88]  =  7'b1110000;     //88pi/512
   cos[88]  =  7'b0011011;     //88pi/512
   sin[89]  =  7'b1101111;     //89pi/512
   cos[89]  =  7'b0011011;     //89pi/512
   sin[90]  =  7'b1101111;     //90pi/512
   cos[90]  =  7'b0011011;     //90pi/512
   sin[91]  =  7'b1101111;     //91pi/512
   cos[91]  =  7'b0011011;     //91pi/512
   sin[92]  =  7'b1101111;     //92pi/512
   cos[92]  =  7'b0011011;     //92pi/512
   sin[93]  =  7'b1101111;     //93pi/512
   cos[93]  =  7'b0011010;     //93pi/512
   sin[94]  =  7'b1101111;     //94pi/512
   cos[94]  =  7'b0011010;     //94pi/512
   sin[95]  =  7'b1101110;     //95pi/512
   cos[95]  =  7'b0011010;     //95pi/512
   sin[96]  =  7'b1101110;     //96pi/512
   cos[96]  =  7'b0011010;     //96pi/512
   sin[97]  =  7'b1101110;     //97pi/512
   cos[97]  =  7'b0011010;     //97pi/512
   sin[98]  =  7'b1101110;     //98pi/512
   cos[98]  =  7'b0011010;     //98pi/512
   sin[99]  =  7'b1101110;     //99pi/512
   cos[99]  =  7'b0011010;     //99pi/512
   sin[100]  =  7'b1101110;     //100pi/512
   cos[100]  =  7'b0011010;     //100pi/512
   sin[101]  =  7'b1101101;     //101pi/512
   cos[101]  =  7'b0011010;     //101pi/512
   sin[102]  =  7'b1101101;     //102pi/512
   cos[102]  =  7'b0011001;     //102pi/512
   sin[103]  =  7'b1101101;     //103pi/512
   cos[103]  =  7'b0011001;     //103pi/512
   sin[104]  =  7'b1101101;     //104pi/512
   cos[104]  =  7'b0011001;     //104pi/512
   sin[105]  =  7'b1101101;     //105pi/512
   cos[105]  =  7'b0011001;     //105pi/512
   sin[106]  =  7'b1101101;     //106pi/512
   cos[106]  =  7'b0011001;     //106pi/512
   sin[107]  =  7'b1101100;     //107pi/512
   cos[107]  =  7'b0011001;     //107pi/512
   sin[108]  =  7'b1101100;     //108pi/512
   cos[108]  =  7'b0011001;     //108pi/512
   sin[109]  =  7'b1101100;     //109pi/512
   cos[109]  =  7'b0011001;     //109pi/512
   sin[110]  =  7'b1101100;     //110pi/512
   cos[110]  =  7'b0011000;     //110pi/512
   sin[111]  =  7'b1101100;     //111pi/512
   cos[111]  =  7'b0011000;     //111pi/512
   sin[112]  =  7'b1101100;     //112pi/512
   cos[112]  =  7'b0011000;     //112pi/512
   sin[113]  =  7'b1101100;     //113pi/512
   cos[113]  =  7'b0011000;     //113pi/512
   sin[114]  =  7'b1101011;     //114pi/512
   cos[114]  =  7'b0011000;     //114pi/512
   sin[115]  =  7'b1101011;     //115pi/512
   cos[115]  =  7'b0011000;     //115pi/512
   sin[116]  =  7'b1101011;     //116pi/512
   cos[116]  =  7'b0011000;     //116pi/512
   sin[117]  =  7'b1101011;     //117pi/512
   cos[117]  =  7'b0011000;     //117pi/512
   sin[118]  =  7'b1101011;     //118pi/512
   cos[118]  =  7'b0010111;     //118pi/512
   sin[119]  =  7'b1101011;     //119pi/512
   cos[119]  =  7'b0010111;     //119pi/512
   sin[120]  =  7'b1101011;     //120pi/512
   cos[120]  =  7'b0010111;     //120pi/512
   sin[121]  =  7'b1101010;     //121pi/512
   cos[121]  =  7'b0010111;     //121pi/512
   sin[122]  =  7'b1101010;     //122pi/512
   cos[122]  =  7'b0010111;     //122pi/512
   sin[123]  =  7'b1101010;     //123pi/512
   cos[123]  =  7'b0010111;     //123pi/512
   sin[124]  =  7'b1101010;     //124pi/512
   cos[124]  =  7'b0010111;     //124pi/512
   sin[125]  =  7'b1101010;     //125pi/512
   cos[125]  =  7'b0010111;     //125pi/512
   sin[126]  =  7'b1101010;     //126pi/512
   cos[126]  =  7'b0010110;     //126pi/512
   sin[127]  =  7'b1101010;     //127pi/512
   cos[127]  =  7'b0010110;     //127pi/512
   sin[128]  =  7'b1101001;     //128pi/512
   cos[128]  =  7'b0010110;     //128pi/512
   sin[129]  =  7'b1101001;     //129pi/512
   cos[129]  =  7'b0010110;     //129pi/512
   sin[130]  =  7'b1101001;     //130pi/512
   cos[130]  =  7'b0010110;     //130pi/512
   sin[131]  =  7'b1101001;     //131pi/512
   cos[131]  =  7'b0010110;     //131pi/512
   sin[132]  =  7'b1101001;     //132pi/512
   cos[132]  =  7'b0010110;     //132pi/512
   sin[133]  =  7'b1101001;     //133pi/512
   cos[133]  =  7'b0010101;     //133pi/512
   sin[134]  =  7'b1101001;     //134pi/512
   cos[134]  =  7'b0010101;     //134pi/512
   sin[135]  =  7'b1101000;     //135pi/512
   cos[135]  =  7'b0010101;     //135pi/512
   sin[136]  =  7'b1101000;     //136pi/512
   cos[136]  =  7'b0010101;     //136pi/512
   sin[137]  =  7'b1101000;     //137pi/512
   cos[137]  =  7'b0010101;     //137pi/512
   sin[138]  =  7'b1101000;     //138pi/512
   cos[138]  =  7'b0010101;     //138pi/512
   sin[139]  =  7'b1101000;     //139pi/512
   cos[139]  =  7'b0010101;     //139pi/512
   sin[140]  =  7'b1101000;     //140pi/512
   cos[140]  =  7'b0010100;     //140pi/512
   sin[141]  =  7'b1101000;     //141pi/512
   cos[141]  =  7'b0010100;     //141pi/512
   sin[142]  =  7'b1101000;     //142pi/512
   cos[142]  =  7'b0010100;     //142pi/512
   sin[143]  =  7'b1100111;     //143pi/512
   cos[143]  =  7'b0010100;     //143pi/512
   sin[144]  =  7'b1100111;     //144pi/512
   cos[144]  =  7'b0010100;     //144pi/512
   sin[145]  =  7'b1100111;     //145pi/512
   cos[145]  =  7'b0010100;     //145pi/512
   sin[146]  =  7'b1100111;     //146pi/512
   cos[146]  =  7'b0010011;     //146pi/512
   sin[147]  =  7'b1100111;     //147pi/512
   cos[147]  =  7'b0010011;     //147pi/512
   sin[148]  =  7'b1100111;     //148pi/512
   cos[148]  =  7'b0010011;     //148pi/512
   sin[149]  =  7'b1100111;     //149pi/512
   cos[149]  =  7'b0010011;     //149pi/512
   sin[150]  =  7'b1100111;     //150pi/512
   cos[150]  =  7'b0010011;     //150pi/512
   sin[151]  =  7'b1100110;     //151pi/512
   cos[151]  =  7'b0010011;     //151pi/512
   sin[152]  =  7'b1100110;     //152pi/512
   cos[152]  =  7'b0010011;     //152pi/512
   sin[153]  =  7'b1100110;     //153pi/512
   cos[153]  =  7'b0010010;     //153pi/512
   sin[154]  =  7'b1100110;     //154pi/512
   cos[154]  =  7'b0010010;     //154pi/512
   sin[155]  =  7'b1100110;     //155pi/512
   cos[155]  =  7'b0010010;     //155pi/512
   sin[156]  =  7'b1100110;     //156pi/512
   cos[156]  =  7'b0010010;     //156pi/512
   sin[157]  =  7'b1100110;     //157pi/512
   cos[157]  =  7'b0010010;     //157pi/512
   sin[158]  =  7'b1100110;     //158pi/512
   cos[158]  =  7'b0010010;     //158pi/512
   sin[159]  =  7'b1100110;     //159pi/512
   cos[159]  =  7'b0010001;     //159pi/512
   sin[160]  =  7'b1100101;     //160pi/512
   cos[160]  =  7'b0010001;     //160pi/512
   sin[161]  =  7'b1100101;     //161pi/512
   cos[161]  =  7'b0010001;     //161pi/512
   sin[162]  =  7'b1100101;     //162pi/512
   cos[162]  =  7'b0010001;     //162pi/512
   sin[163]  =  7'b1100101;     //163pi/512
   cos[163]  =  7'b0010001;     //163pi/512
   sin[164]  =  7'b1100101;     //164pi/512
   cos[164]  =  7'b0010001;     //164pi/512
   sin[165]  =  7'b1100101;     //165pi/512
   cos[165]  =  7'b0010000;     //165pi/512
   sin[166]  =  7'b1100101;     //166pi/512
   cos[166]  =  7'b0010000;     //166pi/512
   sin[167]  =  7'b1100101;     //167pi/512
   cos[167]  =  7'b0010000;     //167pi/512
   sin[168]  =  7'b1100101;     //168pi/512
   cos[168]  =  7'b0010000;     //168pi/512
   sin[169]  =  7'b1100100;     //169pi/512
   cos[169]  =  7'b0010000;     //169pi/512
   sin[170]  =  7'b1100100;     //170pi/512
   cos[170]  =  7'b0010000;     //170pi/512
   sin[171]  =  7'b1100100;     //171pi/512
   cos[171]  =  7'b0001111;     //171pi/512
   sin[172]  =  7'b1100100;     //172pi/512
   cos[172]  =  7'b0001111;     //172pi/512
   sin[173]  =  7'b1100100;     //173pi/512
   cos[173]  =  7'b0001111;     //173pi/512
   sin[174]  =  7'b1100100;     //174pi/512
   cos[174]  =  7'b0001111;     //174pi/512
   sin[175]  =  7'b1100100;     //175pi/512
   cos[175]  =  7'b0001111;     //175pi/512
   sin[176]  =  7'b1100100;     //176pi/512
   cos[176]  =  7'b0001111;     //176pi/512
   sin[177]  =  7'b1100100;     //177pi/512
   cos[177]  =  7'b0001110;     //177pi/512
   sin[178]  =  7'b1100100;     //178pi/512
   cos[178]  =  7'b0001110;     //178pi/512
   sin[179]  =  7'b1100100;     //179pi/512
   cos[179]  =  7'b0001110;     //179pi/512
   sin[180]  =  7'b1100011;     //180pi/512
   cos[180]  =  7'b0001110;     //180pi/512
   sin[181]  =  7'b1100011;     //181pi/512
   cos[181]  =  7'b0001110;     //181pi/512
   sin[182]  =  7'b1100011;     //182pi/512
   cos[182]  =  7'b0001110;     //182pi/512
   sin[183]  =  7'b1100011;     //183pi/512
   cos[183]  =  7'b0001101;     //183pi/512
   sin[184]  =  7'b1100011;     //184pi/512
   cos[184]  =  7'b0001101;     //184pi/512
   sin[185]  =  7'b1100011;     //185pi/512
   cos[185]  =  7'b0001101;     //185pi/512
   sin[186]  =  7'b1100011;     //186pi/512
   cos[186]  =  7'b0001101;     //186pi/512
   sin[187]  =  7'b1100011;     //187pi/512
   cos[187]  =  7'b0001101;     //187pi/512
   sin[188]  =  7'b1100011;     //188pi/512
   cos[188]  =  7'b0001100;     //188pi/512
   sin[189]  =  7'b1100011;     //189pi/512
   cos[189]  =  7'b0001100;     //189pi/512
   sin[190]  =  7'b1100011;     //190pi/512
   cos[190]  =  7'b0001100;     //190pi/512
   sin[191]  =  7'b1100011;     //191pi/512
   cos[191]  =  7'b0001100;     //191pi/512
   sin[192]  =  7'b1100010;     //192pi/512
   cos[192]  =  7'b0001100;     //192pi/512
   sin[193]  =  7'b1100010;     //193pi/512
   cos[193]  =  7'b0001100;     //193pi/512
   sin[194]  =  7'b1100010;     //194pi/512
   cos[194]  =  7'b0001011;     //194pi/512
   sin[195]  =  7'b1100010;     //195pi/512
   cos[195]  =  7'b0001011;     //195pi/512
   sin[196]  =  7'b1100010;     //196pi/512
   cos[196]  =  7'b0001011;     //196pi/512
   sin[197]  =  7'b1100010;     //197pi/512
   cos[197]  =  7'b0001011;     //197pi/512
   sin[198]  =  7'b1100010;     //198pi/512
   cos[198]  =  7'b0001011;     //198pi/512
   sin[199]  =  7'b1100010;     //199pi/512
   cos[199]  =  7'b0001010;     //199pi/512
   sin[200]  =  7'b1100010;     //200pi/512
   cos[200]  =  7'b0001010;     //200pi/512
   sin[201]  =  7'b1100010;     //201pi/512
   cos[201]  =  7'b0001010;     //201pi/512
   sin[202]  =  7'b1100010;     //202pi/512
   cos[202]  =  7'b0001010;     //202pi/512
   sin[203]  =  7'b1100010;     //203pi/512
   cos[203]  =  7'b0001010;     //203pi/512
   sin[204]  =  7'b1100010;     //204pi/512
   cos[204]  =  7'b0001010;     //204pi/512
   sin[205]  =  7'b1100010;     //205pi/512
   cos[205]  =  7'b0001001;     //205pi/512
   sin[206]  =  7'b1100001;     //206pi/512
   cos[206]  =  7'b0001001;     //206pi/512
   sin[207]  =  7'b1100001;     //207pi/512
   cos[207]  =  7'b0001001;     //207pi/512
   sin[208]  =  7'b1100001;     //208pi/512
   cos[208]  =  7'b0001001;     //208pi/512
   sin[209]  =  7'b1100001;     //209pi/512
   cos[209]  =  7'b0001001;     //209pi/512
   sin[210]  =  7'b1100001;     //210pi/512
   cos[210]  =  7'b0001000;     //210pi/512
   sin[211]  =  7'b1100001;     //211pi/512
   cos[211]  =  7'b0001000;     //211pi/512
   sin[212]  =  7'b1100001;     //212pi/512
   cos[212]  =  7'b0001000;     //212pi/512
   sin[213]  =  7'b1100001;     //213pi/512
   cos[213]  =  7'b0001000;     //213pi/512
   sin[214]  =  7'b1100001;     //214pi/512
   cos[214]  =  7'b0001000;     //214pi/512
   sin[215]  =  7'b1100001;     //215pi/512
   cos[215]  =  7'b0000111;     //215pi/512
   sin[216]  =  7'b1100001;     //216pi/512
   cos[216]  =  7'b0000111;     //216pi/512
   sin[217]  =  7'b1100001;     //217pi/512
   cos[217]  =  7'b0000111;     //217pi/512
   sin[218]  =  7'b1100001;     //218pi/512
   cos[218]  =  7'b0000111;     //218pi/512
   sin[219]  =  7'b1100001;     //219pi/512
   cos[219]  =  7'b0000111;     //219pi/512
   sin[220]  =  7'b1100001;     //220pi/512
   cos[220]  =  7'b0000111;     //220pi/512
   sin[221]  =  7'b1100001;     //221pi/512
   cos[221]  =  7'b0000110;     //221pi/512
   sin[222]  =  7'b1100001;     //222pi/512
   cos[222]  =  7'b0000110;     //222pi/512
   sin[223]  =  7'b1100001;     //223pi/512
   cos[223]  =  7'b0000110;     //223pi/512
   sin[224]  =  7'b1100001;     //224pi/512
   cos[224]  =  7'b0000110;     //224pi/512
   sin[225]  =  7'b1100001;     //225pi/512
   cos[225]  =  7'b0000110;     //225pi/512
   sin[226]  =  7'b1100001;     //226pi/512
   cos[226]  =  7'b0000101;     //226pi/512
   sin[227]  =  7'b1100001;     //227pi/512
   cos[227]  =  7'b0000101;     //227pi/512
   sin[228]  =  7'b1100000;     //228pi/512
   cos[228]  =  7'b0000101;     //228pi/512
   sin[229]  =  7'b1100000;     //229pi/512
   cos[229]  =  7'b0000101;     //229pi/512
   sin[230]  =  7'b1100000;     //230pi/512
   cos[230]  =  7'b0000101;     //230pi/512
   sin[231]  =  7'b1100000;     //231pi/512
   cos[231]  =  7'b0000100;     //231pi/512
   sin[232]  =  7'b1100000;     //232pi/512
   cos[232]  =  7'b0000100;     //232pi/512
   sin[233]  =  7'b1100000;     //233pi/512
   cos[233]  =  7'b0000100;     //233pi/512
   sin[234]  =  7'b1100000;     //234pi/512
   cos[234]  =  7'b0000100;     //234pi/512
   sin[235]  =  7'b1100000;     //235pi/512
   cos[235]  =  7'b0000100;     //235pi/512
   sin[236]  =  7'b1100000;     //236pi/512
   cos[236]  =  7'b0000011;     //236pi/512
   sin[237]  =  7'b1100000;     //237pi/512
   cos[237]  =  7'b0000011;     //237pi/512
   sin[238]  =  7'b1100000;     //238pi/512
   cos[238]  =  7'b0000011;     //238pi/512
   sin[239]  =  7'b1100000;     //239pi/512
   cos[239]  =  7'b0000011;     //239pi/512
   sin[240]  =  7'b1100000;     //240pi/512
   cos[240]  =  7'b0000011;     //240pi/512
   sin[241]  =  7'b1100000;     //241pi/512
   cos[241]  =  7'b0000010;     //241pi/512
   sin[242]  =  7'b1100000;     //242pi/512
   cos[242]  =  7'b0000010;     //242pi/512
   sin[243]  =  7'b1100000;     //243pi/512
   cos[243]  =  7'b0000010;     //243pi/512
   sin[244]  =  7'b1100000;     //244pi/512
   cos[244]  =  7'b0000010;     //244pi/512
   sin[245]  =  7'b1100000;     //245pi/512
   cos[245]  =  7'b0000010;     //245pi/512
   sin[246]  =  7'b1100000;     //246pi/512
   cos[246]  =  7'b0000001;     //246pi/512
   sin[247]  =  7'b1100000;     //247pi/512
   cos[247]  =  7'b0000001;     //247pi/512
   sin[248]  =  7'b1100000;     //248pi/512
   cos[248]  =  7'b0000001;     //248pi/512
   sin[249]  =  7'b1100000;     //249pi/512
   cos[249]  =  7'b0000001;     //249pi/512
   sin[250]  =  7'b1100000;     //250pi/512
   cos[250]  =  7'b0000001;     //250pi/512
   sin[251]  =  7'b1100000;     //251pi/512
   cos[251]  =  7'b0000000;     //251pi/512
   sin[252]  =  7'b1100000;     //252pi/512
   cos[252]  =  7'b0000000;     //252pi/512
   sin[253]  =  7'b1100000;     //253pi/512
   cos[253]  =  7'b0000000;     //253pi/512
   sin[254]  =  7'b1100000;     //254pi/512
   cos[254]  =  7'b0000000;     //254pi/512
   sin[255]  =  7'b1100000;     //255pi/512
   cos[255]  =  7'b0000000;     //255pi/512
   sin[256]  =  7'b1100000;     //256pi/512
   cos[256]  =  7'b0000000;     //256pi/512
   sin[257]  =  7'b1100000;     //257pi/512
   cos[257]  =  7'b0000000;     //257pi/512
   sin[258]  =  7'b1100000;     //258pi/512
   cos[258]  =  7'b0000000;     //258pi/512
   sin[259]  =  7'b1100000;     //259pi/512
   cos[259]  =  7'b1111111;     //259pi/512
   sin[260]  =  7'b1100000;     //260pi/512
   cos[260]  =  7'b1111111;     //260pi/512
   sin[261]  =  7'b1100000;     //261pi/512
   cos[261]  =  7'b1111111;     //261pi/512
   sin[262]  =  7'b1100000;     //262pi/512
   cos[262]  =  7'b1111111;     //262pi/512
   sin[263]  =  7'b1100000;     //263pi/512
   cos[263]  =  7'b1111111;     //263pi/512
   sin[264]  =  7'b1100000;     //264pi/512
   cos[264]  =  7'b1111110;     //264pi/512
   sin[265]  =  7'b1100000;     //265pi/512
   cos[265]  =  7'b1111110;     //265pi/512
   sin[266]  =  7'b1100000;     //266pi/512
   cos[266]  =  7'b1111110;     //266pi/512
   sin[267]  =  7'b1100000;     //267pi/512
   cos[267]  =  7'b1111110;     //267pi/512
   sin[268]  =  7'b1100000;     //268pi/512
   cos[268]  =  7'b1111110;     //268pi/512
   sin[269]  =  7'b1100000;     //269pi/512
   cos[269]  =  7'b1111101;     //269pi/512
   sin[270]  =  7'b1100000;     //270pi/512
   cos[270]  =  7'b1111101;     //270pi/512
   sin[271]  =  7'b1100000;     //271pi/512
   cos[271]  =  7'b1111101;     //271pi/512
   sin[272]  =  7'b1100000;     //272pi/512
   cos[272]  =  7'b1111101;     //272pi/512
   sin[273]  =  7'b1100000;     //273pi/512
   cos[273]  =  7'b1111101;     //273pi/512
   sin[274]  =  7'b1100000;     //274pi/512
   cos[274]  =  7'b1111100;     //274pi/512
   sin[275]  =  7'b1100000;     //275pi/512
   cos[275]  =  7'b1111100;     //275pi/512
   sin[276]  =  7'b1100000;     //276pi/512
   cos[276]  =  7'b1111100;     //276pi/512
   sin[277]  =  7'b1100000;     //277pi/512
   cos[277]  =  7'b1111100;     //277pi/512
   sin[278]  =  7'b1100000;     //278pi/512
   cos[278]  =  7'b1111100;     //278pi/512
   sin[279]  =  7'b1100000;     //279pi/512
   cos[279]  =  7'b1111011;     //279pi/512
   sin[280]  =  7'b1100000;     //280pi/512
   cos[280]  =  7'b1111011;     //280pi/512
   sin[281]  =  7'b1100000;     //281pi/512
   cos[281]  =  7'b1111011;     //281pi/512
   sin[282]  =  7'b1100000;     //282pi/512
   cos[282]  =  7'b1111011;     //282pi/512
   sin[283]  =  7'b1100000;     //283pi/512
   cos[283]  =  7'b1111011;     //283pi/512
   sin[284]  =  7'b1100000;     //284pi/512
   cos[284]  =  7'b1111011;     //284pi/512
   sin[285]  =  7'b1100001;     //285pi/512
   cos[285]  =  7'b1111010;     //285pi/512
   sin[286]  =  7'b1100001;     //286pi/512
   cos[286]  =  7'b1111010;     //286pi/512
   sin[287]  =  7'b1100001;     //287pi/512
   cos[287]  =  7'b1111010;     //287pi/512
   sin[288]  =  7'b1100001;     //288pi/512
   cos[288]  =  7'b1111010;     //288pi/512
   sin[289]  =  7'b1100001;     //289pi/512
   cos[289]  =  7'b1111010;     //289pi/512
   sin[290]  =  7'b1100001;     //290pi/512
   cos[290]  =  7'b1111001;     //290pi/512
   sin[291]  =  7'b1100001;     //291pi/512
   cos[291]  =  7'b1111001;     //291pi/512
   sin[292]  =  7'b1100001;     //292pi/512
   cos[292]  =  7'b1111001;     //292pi/512
   sin[293]  =  7'b1100001;     //293pi/512
   cos[293]  =  7'b1111001;     //293pi/512
   sin[294]  =  7'b1100001;     //294pi/512
   cos[294]  =  7'b1111001;     //294pi/512
   sin[295]  =  7'b1100001;     //295pi/512
   cos[295]  =  7'b1111000;     //295pi/512
   sin[296]  =  7'b1100001;     //296pi/512
   cos[296]  =  7'b1111000;     //296pi/512
   sin[297]  =  7'b1100001;     //297pi/512
   cos[297]  =  7'b1111000;     //297pi/512
   sin[298]  =  7'b1100001;     //298pi/512
   cos[298]  =  7'b1111000;     //298pi/512
   sin[299]  =  7'b1100001;     //299pi/512
   cos[299]  =  7'b1111000;     //299pi/512
   sin[300]  =  7'b1100001;     //300pi/512
   cos[300]  =  7'b1110111;     //300pi/512
   sin[301]  =  7'b1100001;     //301pi/512
   cos[301]  =  7'b1110111;     //301pi/512
   sin[302]  =  7'b1100001;     //302pi/512
   cos[302]  =  7'b1110111;     //302pi/512
   sin[303]  =  7'b1100001;     //303pi/512
   cos[303]  =  7'b1110111;     //303pi/512
   sin[304]  =  7'b1100001;     //304pi/512
   cos[304]  =  7'b1110111;     //304pi/512
   sin[305]  =  7'b1100001;     //305pi/512
   cos[305]  =  7'b1110111;     //305pi/512
   sin[306]  =  7'b1100001;     //306pi/512
   cos[306]  =  7'b1110110;     //306pi/512
   sin[307]  =  7'b1100010;     //307pi/512
   cos[307]  =  7'b1110110;     //307pi/512
   sin[308]  =  7'b1100010;     //308pi/512
   cos[308]  =  7'b1110110;     //308pi/512
   sin[309]  =  7'b1100010;     //309pi/512
   cos[309]  =  7'b1110110;     //309pi/512
   sin[310]  =  7'b1100010;     //310pi/512
   cos[310]  =  7'b1110110;     //310pi/512
   sin[311]  =  7'b1100010;     //311pi/512
   cos[311]  =  7'b1110101;     //311pi/512
   sin[312]  =  7'b1100010;     //312pi/512
   cos[312]  =  7'b1110101;     //312pi/512
   sin[313]  =  7'b1100010;     //313pi/512
   cos[313]  =  7'b1110101;     //313pi/512
   sin[314]  =  7'b1100010;     //314pi/512
   cos[314]  =  7'b1110101;     //314pi/512
   sin[315]  =  7'b1100010;     //315pi/512
   cos[315]  =  7'b1110101;     //315pi/512
   sin[316]  =  7'b1100010;     //316pi/512
   cos[316]  =  7'b1110100;     //316pi/512
   sin[317]  =  7'b1100010;     //317pi/512
   cos[317]  =  7'b1110100;     //317pi/512
   sin[318]  =  7'b1100010;     //318pi/512
   cos[318]  =  7'b1110100;     //318pi/512
   sin[319]  =  7'b1100010;     //319pi/512
   cos[319]  =  7'b1110100;     //319pi/512
   sin[320]  =  7'b1100010;     //320pi/512
   cos[320]  =  7'b1110100;     //320pi/512
   sin[321]  =  7'b1100011;     //321pi/512
   cos[321]  =  7'b1110100;     //321pi/512
   sin[322]  =  7'b1100011;     //322pi/512
   cos[322]  =  7'b1110011;     //322pi/512
   sin[323]  =  7'b1100011;     //323pi/512
   cos[323]  =  7'b1110011;     //323pi/512
   sin[324]  =  7'b1100011;     //324pi/512
   cos[324]  =  7'b1110011;     //324pi/512
   sin[325]  =  7'b1100011;     //325pi/512
   cos[325]  =  7'b1110011;     //325pi/512
   sin[326]  =  7'b1100011;     //326pi/512
   cos[326]  =  7'b1110011;     //326pi/512
   sin[327]  =  7'b1100011;     //327pi/512
   cos[327]  =  7'b1110010;     //327pi/512
   sin[328]  =  7'b1100011;     //328pi/512
   cos[328]  =  7'b1110010;     //328pi/512
   sin[329]  =  7'b1100011;     //329pi/512
   cos[329]  =  7'b1110010;     //329pi/512
   sin[330]  =  7'b1100011;     //330pi/512
   cos[330]  =  7'b1110010;     //330pi/512
   sin[331]  =  7'b1100011;     //331pi/512
   cos[331]  =  7'b1110010;     //331pi/512
   sin[332]  =  7'b1100011;     //332pi/512
   cos[332]  =  7'b1110010;     //332pi/512
   sin[333]  =  7'b1100100;     //333pi/512
   cos[333]  =  7'b1110001;     //333pi/512
   sin[334]  =  7'b1100100;     //334pi/512
   cos[334]  =  7'b1110001;     //334pi/512
   sin[335]  =  7'b1100100;     //335pi/512
   cos[335]  =  7'b1110001;     //335pi/512
   sin[336]  =  7'b1100100;     //336pi/512
   cos[336]  =  7'b1110001;     //336pi/512
   sin[337]  =  7'b1100100;     //337pi/512
   cos[337]  =  7'b1110001;     //337pi/512
   sin[338]  =  7'b1100100;     //338pi/512
   cos[338]  =  7'b1110001;     //338pi/512
   sin[339]  =  7'b1100100;     //339pi/512
   cos[339]  =  7'b1110000;     //339pi/512
   sin[340]  =  7'b1100100;     //340pi/512
   cos[340]  =  7'b1110000;     //340pi/512
   sin[341]  =  7'b1100100;     //341pi/512
   cos[341]  =  7'b1110000;     //341pi/512
   sin[342]  =  7'b1100100;     //342pi/512
   cos[342]  =  7'b1110000;     //342pi/512
   sin[343]  =  7'b1100100;     //343pi/512
   cos[343]  =  7'b1110000;     //343pi/512
   sin[344]  =  7'b1100101;     //344pi/512
   cos[344]  =  7'b1110000;     //344pi/512
   sin[345]  =  7'b1100101;     //345pi/512
   cos[345]  =  7'b1101111;     //345pi/512
   sin[346]  =  7'b1100101;     //346pi/512
   cos[346]  =  7'b1101111;     //346pi/512
   sin[347]  =  7'b1100101;     //347pi/512
   cos[347]  =  7'b1101111;     //347pi/512
   sin[348]  =  7'b1100101;     //348pi/512
   cos[348]  =  7'b1101111;     //348pi/512
   sin[349]  =  7'b1100101;     //349pi/512
   cos[349]  =  7'b1101111;     //349pi/512
   sin[350]  =  7'b1100101;     //350pi/512
   cos[350]  =  7'b1101111;     //350pi/512
   sin[351]  =  7'b1100101;     //351pi/512
   cos[351]  =  7'b1101110;     //351pi/512
   sin[352]  =  7'b1100101;     //352pi/512
   cos[352]  =  7'b1101110;     //352pi/512
   sin[353]  =  7'b1100110;     //353pi/512
   cos[353]  =  7'b1101110;     //353pi/512
   sin[354]  =  7'b1100110;     //354pi/512
   cos[354]  =  7'b1101110;     //354pi/512
   sin[355]  =  7'b1100110;     //355pi/512
   cos[355]  =  7'b1101110;     //355pi/512
   sin[356]  =  7'b1100110;     //356pi/512
   cos[356]  =  7'b1101110;     //356pi/512
   sin[357]  =  7'b1100110;     //357pi/512
   cos[357]  =  7'b1101101;     //357pi/512
   sin[358]  =  7'b1100110;     //358pi/512
   cos[358]  =  7'b1101101;     //358pi/512
   sin[359]  =  7'b1100110;     //359pi/512
   cos[359]  =  7'b1101101;     //359pi/512
   sin[360]  =  7'b1100110;     //360pi/512
   cos[360]  =  7'b1101101;     //360pi/512
   sin[361]  =  7'b1100110;     //361pi/512
   cos[361]  =  7'b1101101;     //361pi/512
   sin[362]  =  7'b1100111;     //362pi/512
   cos[362]  =  7'b1101101;     //362pi/512
   sin[363]  =  7'b1100111;     //363pi/512
   cos[363]  =  7'b1101100;     //363pi/512
   sin[364]  =  7'b1100111;     //364pi/512
   cos[364]  =  7'b1101100;     //364pi/512
   sin[365]  =  7'b1100111;     //365pi/512
   cos[365]  =  7'b1101100;     //365pi/512
   sin[366]  =  7'b1100111;     //366pi/512
   cos[366]  =  7'b1101100;     //366pi/512
   sin[367]  =  7'b1100111;     //367pi/512
   cos[367]  =  7'b1101100;     //367pi/512
   sin[368]  =  7'b1100111;     //368pi/512
   cos[368]  =  7'b1101100;     //368pi/512
   sin[369]  =  7'b1100111;     //369pi/512
   cos[369]  =  7'b1101100;     //369pi/512
   sin[370]  =  7'b1101000;     //370pi/512
   cos[370]  =  7'b1101011;     //370pi/512
   sin[371]  =  7'b1101000;     //371pi/512
   cos[371]  =  7'b1101011;     //371pi/512
   sin[372]  =  7'b1101000;     //372pi/512
   cos[372]  =  7'b1101011;     //372pi/512
   sin[373]  =  7'b1101000;     //373pi/512
   cos[373]  =  7'b1101011;     //373pi/512
   sin[374]  =  7'b1101000;     //374pi/512
   cos[374]  =  7'b1101011;     //374pi/512
   sin[375]  =  7'b1101000;     //375pi/512
   cos[375]  =  7'b1101011;     //375pi/512
   sin[376]  =  7'b1101000;     //376pi/512
   cos[376]  =  7'b1101011;     //376pi/512
   sin[377]  =  7'b1101000;     //377pi/512
   cos[377]  =  7'b1101010;     //377pi/512
   sin[378]  =  7'b1101001;     //378pi/512
   cos[378]  =  7'b1101010;     //378pi/512
   sin[379]  =  7'b1101001;     //379pi/512
   cos[379]  =  7'b1101010;     //379pi/512
   sin[380]  =  7'b1101001;     //380pi/512
   cos[380]  =  7'b1101010;     //380pi/512
   sin[381]  =  7'b1101001;     //381pi/512
   cos[381]  =  7'b1101010;     //381pi/512
   sin[382]  =  7'b1101001;     //382pi/512
   cos[382]  =  7'b1101010;     //382pi/512
   sin[383]  =  7'b1101001;     //383pi/512
   cos[383]  =  7'b1101010;     //383pi/512
   sin[384]  =  7'b1101001;     //384pi/512
   cos[384]  =  7'b1101001;     //384pi/512
   sin[385]  =  7'b1101010;     //385pi/512
   cos[385]  =  7'b1101001;     //385pi/512
   sin[386]  =  7'b1101010;     //386pi/512
   cos[386]  =  7'b1101001;     //386pi/512
   sin[387]  =  7'b1101010;     //387pi/512
   cos[387]  =  7'b1101001;     //387pi/512
   sin[388]  =  7'b1101010;     //388pi/512
   cos[388]  =  7'b1101001;     //388pi/512
   sin[389]  =  7'b1101010;     //389pi/512
   cos[389]  =  7'b1101001;     //389pi/512
   sin[390]  =  7'b1101010;     //390pi/512
   cos[390]  =  7'b1101001;     //390pi/512
   sin[391]  =  7'b1101010;     //391pi/512
   cos[391]  =  7'b1101000;     //391pi/512
   sin[392]  =  7'b1101011;     //392pi/512
   cos[392]  =  7'b1101000;     //392pi/512
   sin[393]  =  7'b1101011;     //393pi/512
   cos[393]  =  7'b1101000;     //393pi/512
   sin[394]  =  7'b1101011;     //394pi/512
   cos[394]  =  7'b1101000;     //394pi/512
   sin[395]  =  7'b1101011;     //395pi/512
   cos[395]  =  7'b1101000;     //395pi/512
   sin[396]  =  7'b1101011;     //396pi/512
   cos[396]  =  7'b1101000;     //396pi/512
   sin[397]  =  7'b1101011;     //397pi/512
   cos[397]  =  7'b1101000;     //397pi/512
   sin[398]  =  7'b1101011;     //398pi/512
   cos[398]  =  7'b1101000;     //398pi/512
   sin[399]  =  7'b1101100;     //399pi/512
   cos[399]  =  7'b1100111;     //399pi/512
   sin[400]  =  7'b1101100;     //400pi/512
   cos[400]  =  7'b1100111;     //400pi/512
   sin[401]  =  7'b1101100;     //401pi/512
   cos[401]  =  7'b1100111;     //401pi/512
   sin[402]  =  7'b1101100;     //402pi/512
   cos[402]  =  7'b1100111;     //402pi/512
   sin[403]  =  7'b1101100;     //403pi/512
   cos[403]  =  7'b1100111;     //403pi/512
   sin[404]  =  7'b1101100;     //404pi/512
   cos[404]  =  7'b1100111;     //404pi/512
   sin[405]  =  7'b1101100;     //405pi/512
   cos[405]  =  7'b1100111;     //405pi/512
   sin[406]  =  7'b1101101;     //406pi/512
   cos[406]  =  7'b1100111;     //406pi/512
   sin[407]  =  7'b1101101;     //407pi/512
   cos[407]  =  7'b1100110;     //407pi/512
   sin[408]  =  7'b1101101;     //408pi/512
   cos[408]  =  7'b1100110;     //408pi/512
   sin[409]  =  7'b1101101;     //409pi/512
   cos[409]  =  7'b1100110;     //409pi/512
   sin[410]  =  7'b1101101;     //410pi/512
   cos[410]  =  7'b1100110;     //410pi/512
   sin[411]  =  7'b1101101;     //411pi/512
   cos[411]  =  7'b1100110;     //411pi/512
   sin[412]  =  7'b1101110;     //412pi/512
   cos[412]  =  7'b1100110;     //412pi/512
   sin[413]  =  7'b1101110;     //413pi/512
   cos[413]  =  7'b1100110;     //413pi/512
   sin[414]  =  7'b1101110;     //414pi/512
   cos[414]  =  7'b1100110;     //414pi/512
   sin[415]  =  7'b1101110;     //415pi/512
   cos[415]  =  7'b1100110;     //415pi/512
   sin[416]  =  7'b1101110;     //416pi/512
   cos[416]  =  7'b1100101;     //416pi/512
   sin[417]  =  7'b1101110;     //417pi/512
   cos[417]  =  7'b1100101;     //417pi/512
   sin[418]  =  7'b1101111;     //418pi/512
   cos[418]  =  7'b1100101;     //418pi/512
   sin[419]  =  7'b1101111;     //419pi/512
   cos[419]  =  7'b1100101;     //419pi/512
   sin[420]  =  7'b1101111;     //420pi/512
   cos[420]  =  7'b1100101;     //420pi/512
   sin[421]  =  7'b1101111;     //421pi/512
   cos[421]  =  7'b1100101;     //421pi/512
   sin[422]  =  7'b1101111;     //422pi/512
   cos[422]  =  7'b1100101;     //422pi/512
   sin[423]  =  7'b1101111;     //423pi/512
   cos[423]  =  7'b1100101;     //423pi/512
   sin[424]  =  7'b1110000;     //424pi/512
   cos[424]  =  7'b1100101;     //424pi/512
   sin[425]  =  7'b1110000;     //425pi/512
   cos[425]  =  7'b1100100;     //425pi/512
   sin[426]  =  7'b1110000;     //426pi/512
   cos[426]  =  7'b1100100;     //426pi/512
   sin[427]  =  7'b1110000;     //427pi/512
   cos[427]  =  7'b1100100;     //427pi/512
   sin[428]  =  7'b1110000;     //428pi/512
   cos[428]  =  7'b1100100;     //428pi/512
   sin[429]  =  7'b1110000;     //429pi/512
   cos[429]  =  7'b1100100;     //429pi/512
   sin[430]  =  7'b1110001;     //430pi/512
   cos[430]  =  7'b1100100;     //430pi/512
   sin[431]  =  7'b1110001;     //431pi/512
   cos[431]  =  7'b1100100;     //431pi/512
   sin[432]  =  7'b1110001;     //432pi/512
   cos[432]  =  7'b1100100;     //432pi/512
   sin[433]  =  7'b1110001;     //433pi/512
   cos[433]  =  7'b1100100;     //433pi/512
   sin[434]  =  7'b1110001;     //434pi/512
   cos[434]  =  7'b1100100;     //434pi/512
   sin[435]  =  7'b1110001;     //435pi/512
   cos[435]  =  7'b1100100;     //435pi/512
   sin[436]  =  7'b1110010;     //436pi/512
   cos[436]  =  7'b1100011;     //436pi/512
   sin[437]  =  7'b1110010;     //437pi/512
   cos[437]  =  7'b1100011;     //437pi/512
   sin[438]  =  7'b1110010;     //438pi/512
   cos[438]  =  7'b1100011;     //438pi/512
   sin[439]  =  7'b1110010;     //439pi/512
   cos[439]  =  7'b1100011;     //439pi/512
   sin[440]  =  7'b1110010;     //440pi/512
   cos[440]  =  7'b1100011;     //440pi/512
   sin[441]  =  7'b1110010;     //441pi/512
   cos[441]  =  7'b1100011;     //441pi/512
   sin[442]  =  7'b1110011;     //442pi/512
   cos[442]  =  7'b1100011;     //442pi/512
   sin[443]  =  7'b1110011;     //443pi/512
   cos[443]  =  7'b1100011;     //443pi/512
   sin[444]  =  7'b1110011;     //444pi/512
   cos[444]  =  7'b1100011;     //444pi/512
   sin[445]  =  7'b1110011;     //445pi/512
   cos[445]  =  7'b1100011;     //445pi/512
   sin[446]  =  7'b1110011;     //446pi/512
   cos[446]  =  7'b1100011;     //446pi/512
   sin[447]  =  7'b1110100;     //447pi/512
   cos[447]  =  7'b1100011;     //447pi/512
   sin[448]  =  7'b1110100;     //448pi/512
   cos[448]  =  7'b1100010;     //448pi/512
   sin[449]  =  7'b1110100;     //449pi/512
   cos[449]  =  7'b1100010;     //449pi/512
   sin[450]  =  7'b1110100;     //450pi/512
   cos[450]  =  7'b1100010;     //450pi/512
   sin[451]  =  7'b1110100;     //451pi/512
   cos[451]  =  7'b1100010;     //451pi/512
   sin[452]  =  7'b1110100;     //452pi/512
   cos[452]  =  7'b1100010;     //452pi/512
   sin[453]  =  7'b1110101;     //453pi/512
   cos[453]  =  7'b1100010;     //453pi/512
   sin[454]  =  7'b1110101;     //454pi/512
   cos[454]  =  7'b1100010;     //454pi/512
   sin[455]  =  7'b1110101;     //455pi/512
   cos[455]  =  7'b1100010;     //455pi/512
   sin[456]  =  7'b1110101;     //456pi/512
   cos[456]  =  7'b1100010;     //456pi/512
   sin[457]  =  7'b1110101;     //457pi/512
   cos[457]  =  7'b1100010;     //457pi/512
   sin[458]  =  7'b1110110;     //458pi/512
   cos[458]  =  7'b1100010;     //458pi/512
   sin[459]  =  7'b1110110;     //459pi/512
   cos[459]  =  7'b1100010;     //459pi/512
   sin[460]  =  7'b1110110;     //460pi/512
   cos[460]  =  7'b1100010;     //460pi/512
   sin[461]  =  7'b1110110;     //461pi/512
   cos[461]  =  7'b1100010;     //461pi/512
   sin[462]  =  7'b1110110;     //462pi/512
   cos[462]  =  7'b1100001;     //462pi/512
   sin[463]  =  7'b1110111;     //463pi/512
   cos[463]  =  7'b1100001;     //463pi/512
   sin[464]  =  7'b1110111;     //464pi/512
   cos[464]  =  7'b1100001;     //464pi/512
   sin[465]  =  7'b1110111;     //465pi/512
   cos[465]  =  7'b1100001;     //465pi/512
   sin[466]  =  7'b1110111;     //466pi/512
   cos[466]  =  7'b1100001;     //466pi/512
   sin[467]  =  7'b1110111;     //467pi/512
   cos[467]  =  7'b1100001;     //467pi/512
   sin[468]  =  7'b1110111;     //468pi/512
   cos[468]  =  7'b1100001;     //468pi/512
   sin[469]  =  7'b1111000;     //469pi/512
   cos[469]  =  7'b1100001;     //469pi/512
   sin[470]  =  7'b1111000;     //470pi/512
   cos[470]  =  7'b1100001;     //470pi/512
   sin[471]  =  7'b1111000;     //471pi/512
   cos[471]  =  7'b1100001;     //471pi/512
   sin[472]  =  7'b1111000;     //472pi/512
   cos[472]  =  7'b1100001;     //472pi/512
   sin[473]  =  7'b1111000;     //473pi/512
   cos[473]  =  7'b1100001;     //473pi/512
   sin[474]  =  7'b1111001;     //474pi/512
   cos[474]  =  7'b1100001;     //474pi/512
   sin[475]  =  7'b1111001;     //475pi/512
   cos[475]  =  7'b1100001;     //475pi/512
   sin[476]  =  7'b1111001;     //476pi/512
   cos[476]  =  7'b1100001;     //476pi/512
   sin[477]  =  7'b1111001;     //477pi/512
   cos[477]  =  7'b1100001;     //477pi/512
   sin[478]  =  7'b1111001;     //478pi/512
   cos[478]  =  7'b1100001;     //478pi/512
   sin[479]  =  7'b1111010;     //479pi/512
   cos[479]  =  7'b1100001;     //479pi/512
   sin[480]  =  7'b1111010;     //480pi/512
   cos[480]  =  7'b1100001;     //480pi/512
   sin[481]  =  7'b1111010;     //481pi/512
   cos[481]  =  7'b1100001;     //481pi/512
   sin[482]  =  7'b1111010;     //482pi/512
   cos[482]  =  7'b1100001;     //482pi/512
   sin[483]  =  7'b1111010;     //483pi/512
   cos[483]  =  7'b1100001;     //483pi/512
   sin[484]  =  7'b1111011;     //484pi/512
   cos[484]  =  7'b1100000;     //484pi/512
   sin[485]  =  7'b1111011;     //485pi/512
   cos[485]  =  7'b1100000;     //485pi/512
   sin[486]  =  7'b1111011;     //486pi/512
   cos[486]  =  7'b1100000;     //486pi/512
   sin[487]  =  7'b1111011;     //487pi/512
   cos[487]  =  7'b1100000;     //487pi/512
   sin[488]  =  7'b1111011;     //488pi/512
   cos[488]  =  7'b1100000;     //488pi/512
   sin[489]  =  7'b1111011;     //489pi/512
   cos[489]  =  7'b1100000;     //489pi/512
   sin[490]  =  7'b1111100;     //490pi/512
   cos[490]  =  7'b1100000;     //490pi/512
   sin[491]  =  7'b1111100;     //491pi/512
   cos[491]  =  7'b1100000;     //491pi/512
   sin[492]  =  7'b1111100;     //492pi/512
   cos[492]  =  7'b1100000;     //492pi/512
   sin[493]  =  7'b1111100;     //493pi/512
   cos[493]  =  7'b1100000;     //493pi/512
   sin[494]  =  7'b1111100;     //494pi/512
   cos[494]  =  7'b1100000;     //494pi/512
   sin[495]  =  7'b1111101;     //495pi/512
   cos[495]  =  7'b1100000;     //495pi/512
   sin[496]  =  7'b1111101;     //496pi/512
   cos[496]  =  7'b1100000;     //496pi/512
   sin[497]  =  7'b1111101;     //497pi/512
   cos[497]  =  7'b1100000;     //497pi/512
   sin[498]  =  7'b1111101;     //498pi/512
   cos[498]  =  7'b1100000;     //498pi/512
   sin[499]  =  7'b1111101;     //499pi/512
   cos[499]  =  7'b1100000;     //499pi/512
   sin[500]  =  7'b1111110;     //500pi/512
   cos[500]  =  7'b1100000;     //500pi/512
   sin[501]  =  7'b1111110;     //501pi/512
   cos[501]  =  7'b1100000;     //501pi/512
   sin[502]  =  7'b1111110;     //502pi/512
   cos[502]  =  7'b1100000;     //502pi/512
   sin[503]  =  7'b1111110;     //503pi/512
   cos[503]  =  7'b1100000;     //503pi/512
   sin[504]  =  7'b1111110;     //504pi/512
   cos[504]  =  7'b1100000;     //504pi/512
   sin[505]  =  7'b1111111;     //505pi/512
   cos[505]  =  7'b1100000;     //505pi/512
   sin[506]  =  7'b1111111;     //506pi/512
   cos[506]  =  7'b1100000;     //506pi/512
   sin[507]  =  7'b1111111;     //507pi/512
   cos[507]  =  7'b1100000;     //507pi/512
   sin[508]  =  7'b1111111;     //508pi/512
   cos[508]  =  7'b1100000;     //508pi/512
   sin[509]  =  7'b1111111;     //509pi/512
   cos[509]  =  7'b1100000;     //509pi/512
   sin[510]  =  7'b0000000;     //510pi/512
   cos[510]  =  7'b1100000;     //510pi/512
   sin[511]  =  7'b0000000;     //511pi/512
   cos[511]  =  7'b1100000;     //511pi/512

  ////////////////////////////////////////////////////////
     m_sin[0]  =  7'b0000000;     //0pi/512
   m_cos[0]  =  7'b0100000;     //0pi/512
   m_sin[1]  =  7'b0000000;     //1pi/512
   m_cos[1]  =  7'b0011111;     //1pi/512
   m_sin[2]  =  7'b0000000;     //2pi/512
   m_cos[2]  =  7'b0011111;     //2pi/512
   m_sin[3]  =  7'b0000000;     //3pi/512
   m_cos[3]  =  7'b0011111;     //3pi/512
   m_sin[4]  =  7'b1111111;     //4pi/512
   m_cos[4]  =  7'b0011111;     //4pi/512
   m_sin[5]  =  7'b1111111;     //5pi/512
   m_cos[5]  =  7'b0011111;     //5pi/512
   m_sin[6]  =  7'b1111111;     //6pi/512
   m_cos[6]  =  7'b0011111;     //6pi/512
   m_sin[7]  =  7'b1111111;     //7pi/512
   m_cos[7]  =  7'b0011111;     //7pi/512
   m_sin[8]  =  7'b1111111;     //8pi/512
   m_cos[8]  =  7'b0011111;     //8pi/512
   m_sin[9]  =  7'b1111111;     //9pi/512
   m_cos[9]  =  7'b0011111;     //9pi/512
   m_sin[10]  =  7'b1111110;     //10pi/512
   m_cos[10]  =  7'b0011111;     //10pi/512
   m_sin[11]  =  7'b1111110;     //11pi/512
   m_cos[11]  =  7'b0011111;     //11pi/512
   m_sin[12]  =  7'b1111110;     //12pi/512
   m_cos[12]  =  7'b0011111;     //12pi/512
   m_sin[13]  =  7'b1111110;     //13pi/512
   m_cos[13]  =  7'b0011111;     //13pi/512
   m_sin[14]  =  7'b1111110;     //14pi/512
   m_cos[14]  =  7'b0011111;     //14pi/512
   m_sin[15]  =  7'b1111110;     //15pi/512
   m_cos[15]  =  7'b0011111;     //15pi/512
   m_sin[16]  =  7'b1111101;     //16pi/512
   m_cos[16]  =  7'b0011111;     //16pi/512
   m_sin[17]  =  7'b1111101;     //17pi/512
   m_cos[17]  =  7'b0011111;     //17pi/512
   m_sin[18]  =  7'b1111101;     //18pi/512
   m_cos[18]  =  7'b0011111;     //18pi/512
   m_sin[19]  =  7'b1111101;     //19pi/512
   m_cos[19]  =  7'b0011111;     //19pi/512
   m_sin[20]  =  7'b1111101;     //20pi/512
   m_cos[20]  =  7'b0011111;     //20pi/512
   m_sin[21]  =  7'b1111101;     //21pi/512
   m_cos[21]  =  7'b0011111;     //21pi/512
   m_sin[22]  =  7'b1111101;     //22pi/512
   m_cos[22]  =  7'b0011111;     //22pi/512
   m_sin[23]  =  7'b1111100;     //23pi/512
   m_cos[23]  =  7'b0011111;     //23pi/512
   m_sin[24]  =  7'b1111100;     //24pi/512
   m_cos[24]  =  7'b0011111;     //24pi/512
   m_sin[25]  =  7'b1111100;     //25pi/512
   m_cos[25]  =  7'b0011111;     //25pi/512
   m_sin[26]  =  7'b1111100;     //26pi/512
   m_cos[26]  =  7'b0011111;     //26pi/512
   m_sin[27]  =  7'b1111100;     //27pi/512
   m_cos[27]  =  7'b0011111;     //27pi/512
   m_sin[28]  =  7'b1111100;     //28pi/512
   m_cos[28]  =  7'b0011111;     //28pi/512
   m_sin[29]  =  7'b1111011;     //29pi/512
   m_cos[29]  =  7'b0011111;     //29pi/512
   m_sin[30]  =  7'b1111011;     //30pi/512
   m_cos[30]  =  7'b0011111;     //30pi/512
   m_sin[31]  =  7'b1111011;     //31pi/512
   m_cos[31]  =  7'b0011111;     //31pi/512
   m_sin[32]  =  7'b1111011;     //32pi/512
   m_cos[32]  =  7'b0011111;     //32pi/512
   m_sin[33]  =  7'b1111011;     //33pi/512
   m_cos[33]  =  7'b0011111;     //33pi/512
   m_sin[34]  =  7'b1111011;     //34pi/512
   m_cos[34]  =  7'b0011111;     //34pi/512
   m_sin[35]  =  7'b1111011;     //35pi/512
   m_cos[35]  =  7'b0011111;     //35pi/512
   m_sin[36]  =  7'b1111010;     //36pi/512
   m_cos[36]  =  7'b0011111;     //36pi/512
   m_sin[37]  =  7'b1111010;     //37pi/512
   m_cos[37]  =  7'b0011111;     //37pi/512
   m_sin[38]  =  7'b1111010;     //38pi/512
   m_cos[38]  =  7'b0011111;     //38pi/512
   m_sin[39]  =  7'b1111010;     //39pi/512
   m_cos[39]  =  7'b0011111;     //39pi/512
   m_sin[40]  =  7'b1111010;     //40pi/512
   m_cos[40]  =  7'b0011111;     //40pi/512
   m_sin[41]  =  7'b1111010;     //41pi/512
   m_cos[41]  =  7'b0011111;     //41pi/512
   m_sin[42]  =  7'b1111001;     //42pi/512
   m_cos[42]  =  7'b0011111;     //42pi/512
   m_sin[43]  =  7'b1111001;     //43pi/512
   m_cos[43]  =  7'b0011111;     //43pi/512
   m_sin[44]  =  7'b1111001;     //44pi/512
   m_cos[44]  =  7'b0011111;     //44pi/512
   m_sin[45]  =  7'b1111001;     //45pi/512
   m_cos[45]  =  7'b0011111;     //45pi/512
   m_sin[46]  =  7'b1111001;     //46pi/512
   m_cos[46]  =  7'b0011111;     //46pi/512
   m_sin[47]  =  7'b1111001;     //47pi/512
   m_cos[47]  =  7'b0011111;     //47pi/512
   m_sin[48]  =  7'b1111001;     //48pi/512
   m_cos[48]  =  7'b0011111;     //48pi/512
   m_sin[49]  =  7'b1111000;     //49pi/512
   m_cos[49]  =  7'b0011111;     //49pi/512
   m_sin[50]  =  7'b1111000;     //50pi/512
   m_cos[50]  =  7'b0011111;     //50pi/512
   m_sin[51]  =  7'b1111000;     //51pi/512
   m_cos[51]  =  7'b0011111;     //51pi/512
   m_sin[52]  =  7'b1111000;     //52pi/512
   m_cos[52]  =  7'b0011110;     //52pi/512
   m_sin[53]  =  7'b1111000;     //53pi/512
   m_cos[53]  =  7'b0011110;     //53pi/512
   m_sin[54]  =  7'b1111000;     //54pi/512
   m_cos[54]  =  7'b0011110;     //54pi/512
   m_sin[55]  =  7'b1110111;     //55pi/512
   m_cos[55]  =  7'b0011110;     //55pi/512
   m_sin[56]  =  7'b1110111;     //56pi/512
   m_cos[56]  =  7'b0011110;     //56pi/512
   m_sin[57]  =  7'b1110111;     //57pi/512
   m_cos[57]  =  7'b0011110;     //57pi/512
   m_sin[58]  =  7'b1110111;     //58pi/512
   m_cos[58]  =  7'b0011110;     //58pi/512
   m_sin[59]  =  7'b1110111;     //59pi/512
   m_cos[59]  =  7'b0011110;     //59pi/512
   m_sin[60]  =  7'b1110111;     //60pi/512
   m_cos[60]  =  7'b0011110;     //60pi/512
   m_sin[61]  =  7'b1110111;     //61pi/512
   m_cos[61]  =  7'b0011110;     //61pi/512
   m_sin[62]  =  7'b1110110;     //62pi/512
   m_cos[62]  =  7'b0011110;     //62pi/512
   m_sin[63]  =  7'b1110110;     //63pi/512
   m_cos[63]  =  7'b0011110;     //63pi/512
   m_sin[64]  =  7'b1110110;     //64pi/512
   m_cos[64]  =  7'b0011110;     //64pi/512
   m_sin[65]  =  7'b1110110;     //65pi/512
   m_cos[65]  =  7'b0011110;     //65pi/512
   m_sin[66]  =  7'b1110110;     //66pi/512
   m_cos[66]  =  7'b0011110;     //66pi/512
   m_sin[67]  =  7'b1110110;     //67pi/512
   m_cos[67]  =  7'b0011110;     //67pi/512
   m_sin[68]  =  7'b1110110;     //68pi/512
   m_cos[68]  =  7'b0011110;     //68pi/512
   m_sin[69]  =  7'b1110101;     //69pi/512
   m_cos[69]  =  7'b0011110;     //69pi/512
   m_sin[70]  =  7'b1110101;     //70pi/512
   m_cos[70]  =  7'b0011110;     //70pi/512
   m_sin[71]  =  7'b1110101;     //71pi/512
   m_cos[71]  =  7'b0011110;     //71pi/512
   m_sin[72]  =  7'b1110101;     //72pi/512
   m_cos[72]  =  7'b0011110;     //72pi/512
   m_sin[73]  =  7'b1110101;     //73pi/512
   m_cos[73]  =  7'b0011101;     //73pi/512
   m_sin[74]  =  7'b1110101;     //74pi/512
   m_cos[74]  =  7'b0011101;     //74pi/512
   m_sin[75]  =  7'b1110100;     //75pi/512
   m_cos[75]  =  7'b0011101;     //75pi/512
   m_sin[76]  =  7'b1110100;     //76pi/512
   m_cos[76]  =  7'b0011101;     //76pi/512
   m_sin[77]  =  7'b1110100;     //77pi/512
   m_cos[77]  =  7'b0011101;     //77pi/512
   m_sin[78]  =  7'b1110100;     //78pi/512
   m_cos[78]  =  7'b0011101;     //78pi/512
   m_sin[79]  =  7'b1110100;     //79pi/512
   m_cos[79]  =  7'b0011101;     //79pi/512
   m_sin[80]  =  7'b1110100;     //80pi/512
   m_cos[80]  =  7'b0011101;     //80pi/512
   m_sin[81]  =  7'b1110100;     //81pi/512
   m_cos[81]  =  7'b0011101;     //81pi/512
   m_sin[82]  =  7'b1110011;     //82pi/512
   m_cos[82]  =  7'b0011101;     //82pi/512
   m_sin[83]  =  7'b1110011;     //83pi/512
   m_cos[83]  =  7'b0011101;     //83pi/512
   m_sin[84]  =  7'b1110011;     //84pi/512
   m_cos[84]  =  7'b0011101;     //84pi/512
   m_sin[85]  =  7'b1110011;     //85pi/512
   m_cos[85]  =  7'b0011101;     //85pi/512
   m_sin[86]  =  7'b1110011;     //86pi/512
   m_cos[86]  =  7'b0011101;     //86pi/512
   m_sin[87]  =  7'b1110011;     //87pi/512
   m_cos[87]  =  7'b0011101;     //87pi/512
   m_sin[88]  =  7'b1110011;     //88pi/512
   m_cos[88]  =  7'b0011101;     //88pi/512
   m_sin[89]  =  7'b1110010;     //89pi/512
   m_cos[89]  =  7'b0011100;     //89pi/512
   m_sin[90]  =  7'b1110010;     //90pi/512
   m_cos[90]  =  7'b0011100;     //90pi/512
   m_sin[91]  =  7'b1110010;     //91pi/512
   m_cos[91]  =  7'b0011100;     //91pi/512
   m_sin[92]  =  7'b1110010;     //92pi/512
   m_cos[92]  =  7'b0011100;     //92pi/512
   m_sin[93]  =  7'b1110010;     //93pi/512
   m_cos[93]  =  7'b0011100;     //93pi/512
   m_sin[94]  =  7'b1110010;     //94pi/512
   m_cos[94]  =  7'b0011100;     //94pi/512
   m_sin[95]  =  7'b1110010;     //95pi/512
   m_cos[95]  =  7'b0011100;     //95pi/512
   m_sin[96]  =  7'b1110001;     //96pi/512
   m_cos[96]  =  7'b0011100;     //96pi/512
   m_sin[97]  =  7'b1110001;     //97pi/512
   m_cos[97]  =  7'b0011100;     //97pi/512
   m_sin[98]  =  7'b1110001;     //98pi/512
   m_cos[98]  =  7'b0011100;     //98pi/512
   m_sin[99]  =  7'b1110001;     //99pi/512
   m_cos[99]  =  7'b0011100;     //99pi/512
   m_sin[100]  =  7'b1110001;     //100pi/512
   m_cos[100]  =  7'b0011100;     //100pi/512
   m_sin[101]  =  7'b1110001;     //101pi/512
   m_cos[101]  =  7'b0011100;     //101pi/512
   m_sin[102]  =  7'b1110001;     //102pi/512
   m_cos[102]  =  7'b0011100;     //102pi/512
   m_sin[103]  =  7'b1110001;     //103pi/512
   m_cos[103]  =  7'b0011011;     //103pi/512
   m_sin[104]  =  7'b1110000;     //104pi/512
   m_cos[104]  =  7'b0011011;     //104pi/512
   m_sin[105]  =  7'b1110000;     //105pi/512
   m_cos[105]  =  7'b0011011;     //105pi/512
   m_sin[106]  =  7'b1110000;     //106pi/512
   m_cos[106]  =  7'b0011011;     //106pi/512
   m_sin[107]  =  7'b1110000;     //107pi/512
   m_cos[107]  =  7'b0011011;     //107pi/512
   m_sin[108]  =  7'b1110000;     //108pi/512
   m_cos[108]  =  7'b0011011;     //108pi/512
   m_sin[109]  =  7'b1110000;     //109pi/512
   m_cos[109]  =  7'b0011011;     //109pi/512
   m_sin[110]  =  7'b1110000;     //110pi/512
   m_cos[110]  =  7'b0011011;     //110pi/512
   m_sin[111]  =  7'b1101111;     //111pi/512
   m_cos[111]  =  7'b0011011;     //111pi/512
   m_sin[112]  =  7'b1101111;     //112pi/512
   m_cos[112]  =  7'b0011011;     //112pi/512
   m_sin[113]  =  7'b1101111;     //113pi/512
   m_cos[113]  =  7'b0011011;     //113pi/512
   m_sin[114]  =  7'b1101111;     //114pi/512
   m_cos[114]  =  7'b0011011;     //114pi/512
   m_sin[115]  =  7'b1101111;     //115pi/512
   m_cos[115]  =  7'b0011011;     //115pi/512
   m_sin[116]  =  7'b1101111;     //116pi/512
   m_cos[116]  =  7'b0011010;     //116pi/512
   m_sin[117]  =  7'b1101111;     //117pi/512
   m_cos[117]  =  7'b0011010;     //117pi/512
   m_sin[118]  =  7'b1101110;     //118pi/512
   m_cos[118]  =  7'b0011010;     //118pi/512
   m_sin[119]  =  7'b1101110;     //119pi/512
   m_cos[119]  =  7'b0011010;     //119pi/512
   m_sin[120]  =  7'b1101110;     //120pi/512
   m_cos[120]  =  7'b0011010;     //120pi/512
   m_sin[121]  =  7'b1101110;     //121pi/512
   m_cos[121]  =  7'b0011010;     //121pi/512
   m_sin[122]  =  7'b1101110;     //122pi/512
   m_cos[122]  =  7'b0011010;     //122pi/512
   m_sin[123]  =  7'b1101110;     //123pi/512
   m_cos[123]  =  7'b0011010;     //123pi/512
   m_sin[124]  =  7'b1101110;     //124pi/512
   m_cos[124]  =  7'b0011010;     //124pi/512
   m_sin[125]  =  7'b1101110;     //125pi/512
   m_cos[125]  =  7'b0011010;     //125pi/512
   m_sin[126]  =  7'b1101101;     //126pi/512
   m_cos[126]  =  7'b0011010;     //126pi/512
   m_sin[127]  =  7'b1101101;     //127pi/512
   m_cos[127]  =  7'b0011001;     //127pi/512
   m_sin[128]  =  7'b1101101;     //128pi/512
   m_cos[128]  =  7'b0011001;     //128pi/512
   m_sin[129]  =  7'b1101101;     //129pi/512
   m_cos[129]  =  7'b0011001;     //129pi/512
   m_sin[130]  =  7'b1101101;     //130pi/512
   m_cos[130]  =  7'b0011001;     //130pi/512
   m_sin[131]  =  7'b1101101;     //131pi/512
   m_cos[131]  =  7'b0011001;     //131pi/512
   m_sin[132]  =  7'b1101101;     //132pi/512
   m_cos[132]  =  7'b0011001;     //132pi/512
   m_sin[133]  =  7'b1101101;     //133pi/512
   m_cos[133]  =  7'b0011001;     //133pi/512
   m_sin[134]  =  7'b1101100;     //134pi/512
   m_cos[134]  =  7'b0011001;     //134pi/512
   m_sin[135]  =  7'b1101100;     //135pi/512
   m_cos[135]  =  7'b0011001;     //135pi/512
   m_sin[136]  =  7'b1101100;     //136pi/512
   m_cos[136]  =  7'b0011001;     //136pi/512
   m_sin[137]  =  7'b1101100;     //137pi/512
   m_cos[137]  =  7'b0011001;     //137pi/512
   m_sin[138]  =  7'b1101100;     //138pi/512
   m_cos[138]  =  7'b0011000;     //138pi/512
   m_sin[139]  =  7'b1101100;     //139pi/512
   m_cos[139]  =  7'b0011000;     //139pi/512
   m_sin[140]  =  7'b1101100;     //140pi/512
   m_cos[140]  =  7'b0011000;     //140pi/512
   m_sin[141]  =  7'b1101100;     //141pi/512
   m_cos[141]  =  7'b0011000;     //141pi/512
   m_sin[142]  =  7'b1101011;     //142pi/512
   m_cos[142]  =  7'b0011000;     //142pi/512
   m_sin[143]  =  7'b1101011;     //143pi/512
   m_cos[143]  =  7'b0011000;     //143pi/512
   m_sin[144]  =  7'b1101011;     //144pi/512
   m_cos[144]  =  7'b0011000;     //144pi/512
   m_sin[145]  =  7'b1101011;     //145pi/512
   m_cos[145]  =  7'b0011000;     //145pi/512
   m_sin[146]  =  7'b1101011;     //146pi/512
   m_cos[146]  =  7'b0011000;     //146pi/512
   m_sin[147]  =  7'b1101011;     //147pi/512
   m_cos[147]  =  7'b0011000;     //147pi/512
   m_sin[148]  =  7'b1101011;     //148pi/512
   m_cos[148]  =  7'b0010111;     //148pi/512
   m_sin[149]  =  7'b1101011;     //149pi/512
   m_cos[149]  =  7'b0010111;     //149pi/512
   m_sin[150]  =  7'b1101011;     //150pi/512
   m_cos[150]  =  7'b0010111;     //150pi/512
   m_sin[151]  =  7'b1101010;     //151pi/512
   m_cos[151]  =  7'b0010111;     //151pi/512
   m_sin[152]  =  7'b1101010;     //152pi/512
   m_cos[152]  =  7'b0010111;     //152pi/512
   m_sin[153]  =  7'b1101010;     //153pi/512
   m_cos[153]  =  7'b0010111;     //153pi/512
   m_sin[154]  =  7'b1101010;     //154pi/512
   m_cos[154]  =  7'b0010111;     //154pi/512
   m_sin[155]  =  7'b1101010;     //155pi/512
   m_cos[155]  =  7'b0010111;     //155pi/512
   m_sin[156]  =  7'b1101010;     //156pi/512
   m_cos[156]  =  7'b0010111;     //156pi/512
   m_sin[157]  =  7'b1101010;     //157pi/512
   m_cos[157]  =  7'b0010110;     //157pi/512
   m_sin[158]  =  7'b1101010;     //158pi/512
   m_cos[158]  =  7'b0010110;     //158pi/512
   m_sin[159]  =  7'b1101001;     //159pi/512
   m_cos[159]  =  7'b0010110;     //159pi/512
   m_sin[160]  =  7'b1101001;     //160pi/512
   m_cos[160]  =  7'b0010110;     //160pi/512
   m_sin[161]  =  7'b1101001;     //161pi/512
   m_cos[161]  =  7'b0010110;     //161pi/512
   m_sin[162]  =  7'b1101001;     //162pi/512
   m_cos[162]  =  7'b0010110;     //162pi/512
   m_sin[163]  =  7'b1101001;     //163pi/512
   m_cos[163]  =  7'b0010110;     //163pi/512
   m_sin[164]  =  7'b1101001;     //164pi/512
   m_cos[164]  =  7'b0010110;     //164pi/512
   m_sin[165]  =  7'b1101001;     //165pi/512
   m_cos[165]  =  7'b0010110;     //165pi/512
   m_sin[166]  =  7'b1101001;     //166pi/512
   m_cos[166]  =  7'b0010101;     //166pi/512
   m_sin[167]  =  7'b1101001;     //167pi/512
   m_cos[167]  =  7'b0010101;     //167pi/512
   m_sin[168]  =  7'b1101001;     //168pi/512
   m_cos[168]  =  7'b0010101;     //168pi/512
   m_sin[169]  =  7'b1101000;     //169pi/512
   m_cos[169]  =  7'b0010101;     //169pi/512
   m_sin[170]  =  7'b1101000;     //170pi/512
   m_cos[170]  =  7'b0010101;     //170pi/512
   m_sin[171]  =  7'b1101000;     //171pi/512
   m_cos[171]  =  7'b0010101;     //171pi/512
   m_sin[172]  =  7'b1101000;     //172pi/512
   m_cos[172]  =  7'b0010101;     //172pi/512
   m_sin[173]  =  7'b1101000;     //173pi/512
   m_cos[173]  =  7'b0010101;     //173pi/512
   m_sin[174]  =  7'b1101000;     //174pi/512
   m_cos[174]  =  7'b0010101;     //174pi/512
   m_sin[175]  =  7'b1101000;     //175pi/512
   m_cos[175]  =  7'b0010100;     //175pi/512
   m_sin[176]  =  7'b1101000;     //176pi/512
   m_cos[176]  =  7'b0010100;     //176pi/512
   m_sin[177]  =  7'b1101000;     //177pi/512
   m_cos[177]  =  7'b0010100;     //177pi/512
   m_sin[178]  =  7'b1100111;     //178pi/512
   m_cos[178]  =  7'b0010100;     //178pi/512
   m_sin[179]  =  7'b1100111;     //179pi/512
   m_cos[179]  =  7'b0010100;     //179pi/512
   m_sin[180]  =  7'b1100111;     //180pi/512
   m_cos[180]  =  7'b0010100;     //180pi/512
   m_sin[181]  =  7'b1100111;     //181pi/512
   m_cos[181]  =  7'b0010100;     //181pi/512
   m_sin[182]  =  7'b1100111;     //182pi/512
   m_cos[182]  =  7'b0010100;     //182pi/512
   m_sin[183]  =  7'b1100111;     //183pi/512
   m_cos[183]  =  7'b0010011;     //183pi/512
   m_sin[184]  =  7'b1100111;     //184pi/512
   m_cos[184]  =  7'b0010011;     //184pi/512
   m_sin[185]  =  7'b1100111;     //185pi/512
   m_cos[185]  =  7'b0010011;     //185pi/512
   m_sin[186]  =  7'b1100111;     //186pi/512
   m_cos[186]  =  7'b0010011;     //186pi/512
   m_sin[187]  =  7'b1100111;     //187pi/512
   m_cos[187]  =  7'b0010011;     //187pi/512
   m_sin[188]  =  7'b1100110;     //188pi/512
   m_cos[188]  =  7'b0010011;     //188pi/512
   m_sin[189]  =  7'b1100110;     //189pi/512
   m_cos[189]  =  7'b0010011;     //189pi/512
   m_sin[190]  =  7'b1100110;     //190pi/512
   m_cos[190]  =  7'b0010011;     //190pi/512
   m_sin[191]  =  7'b1100110;     //191pi/512
   m_cos[191]  =  7'b0010010;     //191pi/512
   m_sin[192]  =  7'b1100110;     //192pi/512
   m_cos[192]  =  7'b0010010;     //192pi/512
   m_sin[193]  =  7'b1100110;     //193pi/512
   m_cos[193]  =  7'b0010010;     //193pi/512
   m_sin[194]  =  7'b1100110;     //194pi/512
   m_cos[194]  =  7'b0010010;     //194pi/512
   m_sin[195]  =  7'b1100110;     //195pi/512
   m_cos[195]  =  7'b0010010;     //195pi/512
   m_sin[196]  =  7'b1100110;     //196pi/512
   m_cos[196]  =  7'b0010010;     //196pi/512
   m_sin[197]  =  7'b1100110;     //197pi/512
   m_cos[197]  =  7'b0010010;     //197pi/512
   m_sin[198]  =  7'b1100110;     //198pi/512
   m_cos[198]  =  7'b0010010;     //198pi/512
   m_sin[199]  =  7'b1100101;     //199pi/512
   m_cos[199]  =  7'b0010001;     //199pi/512
   m_sin[200]  =  7'b1100101;     //200pi/512
   m_cos[200]  =  7'b0010001;     //200pi/512
   m_sin[201]  =  7'b1100101;     //201pi/512
   m_cos[201]  =  7'b0010001;     //201pi/512
   m_sin[202]  =  7'b1100101;     //202pi/512
   m_cos[202]  =  7'b0010001;     //202pi/512
   m_sin[203]  =  7'b1100101;     //203pi/512
   m_cos[203]  =  7'b0010001;     //203pi/512
   m_sin[204]  =  7'b1100101;     //204pi/512
   m_cos[204]  =  7'b0010001;     //204pi/512
   m_sin[205]  =  7'b1100101;     //205pi/512
   m_cos[205]  =  7'b0010001;     //205pi/512
   m_sin[206]  =  7'b1100101;     //206pi/512
   m_cos[206]  =  7'b0010000;     //206pi/512
   m_sin[207]  =  7'b1100101;     //207pi/512
   m_cos[207]  =  7'b0010000;     //207pi/512
   m_sin[208]  =  7'b1100101;     //208pi/512
   m_cos[208]  =  7'b0010000;     //208pi/512
   m_sin[209]  =  7'b1100101;     //209pi/512
   m_cos[209]  =  7'b0010000;     //209pi/512
   m_sin[210]  =  7'b1100101;     //210pi/512
   m_cos[210]  =  7'b0010000;     //210pi/512
   m_sin[211]  =  7'b1100100;     //211pi/512
   m_cos[211]  =  7'b0010000;     //211pi/512
   m_sin[212]  =  7'b1100100;     //212pi/512
   m_cos[212]  =  7'b0010000;     //212pi/512
   m_sin[213]  =  7'b1100100;     //213pi/512
   m_cos[213]  =  7'b0010000;     //213pi/512
   m_sin[214]  =  7'b1100100;     //214pi/512
   m_cos[214]  =  7'b0001111;     //214pi/512
   m_sin[215]  =  7'b1100100;     //215pi/512
   m_cos[215]  =  7'b0001111;     //215pi/512
   m_sin[216]  =  7'b1100100;     //216pi/512
   m_cos[216]  =  7'b0001111;     //216pi/512
   m_sin[217]  =  7'b1100100;     //217pi/512
   m_cos[217]  =  7'b0001111;     //217pi/512
   m_sin[218]  =  7'b1100100;     //218pi/512
   m_cos[218]  =  7'b0001111;     //218pi/512
   m_sin[219]  =  7'b1100100;     //219pi/512
   m_cos[219]  =  7'b0001111;     //219pi/512
   m_sin[220]  =  7'b1100100;     //220pi/512
   m_cos[220]  =  7'b0001111;     //220pi/512
   m_sin[221]  =  7'b1100100;     //221pi/512
   m_cos[221]  =  7'b0001110;     //221pi/512
   m_sin[222]  =  7'b1100100;     //222pi/512
   m_cos[222]  =  7'b0001110;     //222pi/512
   m_sin[223]  =  7'b1100100;     //223pi/512
   m_cos[223]  =  7'b0001110;     //223pi/512
   m_sin[224]  =  7'b1100011;     //224pi/512
   m_cos[224]  =  7'b0001110;     //224pi/512
   m_sin[225]  =  7'b1100011;     //225pi/512
   m_cos[225]  =  7'b0001110;     //225pi/512
   m_sin[226]  =  7'b1100011;     //226pi/512
   m_cos[226]  =  7'b0001110;     //226pi/512
   m_sin[227]  =  7'b1100011;     //227pi/512
   m_cos[227]  =  7'b0001110;     //227pi/512
   m_sin[228]  =  7'b1100011;     //228pi/512
   m_cos[228]  =  7'b0001101;     //228pi/512
   m_sin[229]  =  7'b1100011;     //229pi/512
   m_cos[229]  =  7'b0001101;     //229pi/512
   m_sin[230]  =  7'b1100011;     //230pi/512
   m_cos[230]  =  7'b0001101;     //230pi/512
   m_sin[231]  =  7'b1100011;     //231pi/512
   m_cos[231]  =  7'b0001101;     //231pi/512
   m_sin[232]  =  7'b1100011;     //232pi/512
   m_cos[232]  =  7'b0001101;     //232pi/512
   m_sin[233]  =  7'b1100011;     //233pi/512
   m_cos[233]  =  7'b0001101;     //233pi/512
   m_sin[234]  =  7'b1100011;     //234pi/512
   m_cos[234]  =  7'b0001101;     //234pi/512
   m_sin[235]  =  7'b1100011;     //235pi/512
   m_cos[235]  =  7'b0001100;     //235pi/512
   m_sin[236]  =  7'b1100011;     //236pi/512
   m_cos[236]  =  7'b0001100;     //236pi/512
   m_sin[237]  =  7'b1100011;     //237pi/512
   m_cos[237]  =  7'b0001100;     //237pi/512
   m_sin[238]  =  7'b1100011;     //238pi/512
   m_cos[238]  =  7'b0001100;     //238pi/512
   m_sin[239]  =  7'b1100010;     //239pi/512
   m_cos[239]  =  7'b0001100;     //239pi/512
   m_sin[240]  =  7'b1100010;     //240pi/512
   m_cos[240]  =  7'b0001100;     //240pi/512
   m_sin[241]  =  7'b1100010;     //241pi/512
   m_cos[241]  =  7'b0001100;     //241pi/512
   m_sin[242]  =  7'b1100010;     //242pi/512
   m_cos[242]  =  7'b0001011;     //242pi/512
   m_sin[243]  =  7'b1100010;     //243pi/512
   m_cos[243]  =  7'b0001011;     //243pi/512
   m_sin[244]  =  7'b1100010;     //244pi/512
   m_cos[244]  =  7'b0001011;     //244pi/512
   m_sin[245]  =  7'b1100010;     //245pi/512
   m_cos[245]  =  7'b0001011;     //245pi/512
   m_sin[246]  =  7'b1100010;     //246pi/512
   m_cos[246]  =  7'b0001011;     //246pi/512
   m_sin[247]  =  7'b1100010;     //247pi/512
   m_cos[247]  =  7'b0001011;     //247pi/512
   m_sin[248]  =  7'b1100010;     //248pi/512
   m_cos[248]  =  7'b0001011;     //248pi/512
   m_sin[249]  =  7'b1100010;     //249pi/512
   m_cos[249]  =  7'b0001010;     //249pi/512
   m_sin[250]  =  7'b1100010;     //250pi/512
   m_cos[250]  =  7'b0001010;     //250pi/512
   m_sin[251]  =  7'b1100010;     //251pi/512
   m_cos[251]  =  7'b0001010;     //251pi/512
   m_sin[252]  =  7'b1100010;     //252pi/512
   m_cos[252]  =  7'b0001010;     //252pi/512
   m_sin[253]  =  7'b1100010;     //253pi/512
   m_cos[253]  =  7'b0001010;     //253pi/512
   m_sin[254]  =  7'b1100010;     //254pi/512
   m_cos[254]  =  7'b0001010;     //254pi/512
   m_sin[255]  =  7'b1100010;     //255pi/512
   m_cos[255]  =  7'b0001010;     //255pi/512
   m_sin[256]  =  7'b1100010;     //256pi/512
   m_cos[256]  =  7'b0001001;     //256pi/512
   m_sin[257]  =  7'b1100010;     //257pi/512
   m_cos[257]  =  7'b0001001;     //257pi/512
   m_sin[258]  =  7'b1100001;     //258pi/512
   m_cos[258]  =  7'b0001001;     //258pi/512
   m_sin[259]  =  7'b1100001;     //259pi/512
   m_cos[259]  =  7'b0001001;     //259pi/512
   m_sin[260]  =  7'b1100001;     //260pi/512
   m_cos[260]  =  7'b0001001;     //260pi/512
   m_sin[261]  =  7'b1100001;     //261pi/512
   m_cos[261]  =  7'b0001001;     //261pi/512
   m_sin[262]  =  7'b1100001;     //262pi/512
   m_cos[262]  =  7'b0001000;     //262pi/512
   m_sin[263]  =  7'b1100001;     //263pi/512
   m_cos[263]  =  7'b0001000;     //263pi/512
   m_sin[264]  =  7'b1100001;     //264pi/512
   m_cos[264]  =  7'b0001000;     //264pi/512
   m_sin[265]  =  7'b1100001;     //265pi/512
   m_cos[265]  =  7'b0001000;     //265pi/512
   m_sin[266]  =  7'b1100001;     //266pi/512
   m_cos[266]  =  7'b0001000;     //266pi/512
   m_sin[267]  =  7'b1100001;     //267pi/512
   m_cos[267]  =  7'b0001000;     //267pi/512
   m_sin[268]  =  7'b1100001;     //268pi/512
   m_cos[268]  =  7'b0001000;     //268pi/512
   m_sin[269]  =  7'b1100001;     //269pi/512
   m_cos[269]  =  7'b0000111;     //269pi/512
   m_sin[270]  =  7'b1100001;     //270pi/512
   m_cos[270]  =  7'b0000111;     //270pi/512
   m_sin[271]  =  7'b1100001;     //271pi/512
   m_cos[271]  =  7'b0000111;     //271pi/512
   m_sin[272]  =  7'b1100001;     //272pi/512
   m_cos[272]  =  7'b0000111;     //272pi/512
   m_sin[273]  =  7'b1100001;     //273pi/512
   m_cos[273]  =  7'b0000111;     //273pi/512
   m_sin[274]  =  7'b1100001;     //274pi/512
   m_cos[274]  =  7'b0000111;     //274pi/512
   m_sin[275]  =  7'b1100001;     //275pi/512
   m_cos[275]  =  7'b0000111;     //275pi/512
   m_sin[276]  =  7'b1100001;     //276pi/512
   m_cos[276]  =  7'b0000110;     //276pi/512
   m_sin[277]  =  7'b1100001;     //277pi/512
   m_cos[277]  =  7'b0000110;     //277pi/512
   m_sin[278]  =  7'b1100001;     //278pi/512
   m_cos[278]  =  7'b0000110;     //278pi/512
   m_sin[279]  =  7'b1100001;     //279pi/512
   m_cos[279]  =  7'b0000110;     //279pi/512
   m_sin[280]  =  7'b1100001;     //280pi/512
   m_cos[280]  =  7'b0000110;     //280pi/512
   m_sin[281]  =  7'b1100001;     //281pi/512
   m_cos[281]  =  7'b0000110;     //281pi/512
   m_sin[282]  =  7'b1100001;     //282pi/512
   m_cos[282]  =  7'b0000101;     //282pi/512
   m_sin[283]  =  7'b1100001;     //283pi/512
   m_cos[283]  =  7'b0000101;     //283pi/512
   m_sin[284]  =  7'b1100000;     //284pi/512
   m_cos[284]  =  7'b0000101;     //284pi/512
   m_sin[285]  =  7'b1100000;     //285pi/512
   m_cos[285]  =  7'b0000101;     //285pi/512
   m_sin[286]  =  7'b1100000;     //286pi/512
   m_cos[286]  =  7'b0000101;     //286pi/512
   m_sin[287]  =  7'b1100000;     //287pi/512
   m_cos[287]  =  7'b0000101;     //287pi/512
   m_sin[288]  =  7'b1100000;     //288pi/512
   m_cos[288]  =  7'b0000101;     //288pi/512
   m_sin[289]  =  7'b1100000;     //289pi/512
   m_cos[289]  =  7'b0000100;     //289pi/512
   m_sin[290]  =  7'b1100000;     //290pi/512
   m_cos[290]  =  7'b0000100;     //290pi/512
   m_sin[291]  =  7'b1100000;     //291pi/512
   m_cos[291]  =  7'b0000100;     //291pi/512
   m_sin[292]  =  7'b1100000;     //292pi/512
   m_cos[292]  =  7'b0000100;     //292pi/512
   m_sin[293]  =  7'b1100000;     //293pi/512
   m_cos[293]  =  7'b0000100;     //293pi/512
   m_sin[294]  =  7'b1100000;     //294pi/512
   m_cos[294]  =  7'b0000100;     //294pi/512
   m_sin[295]  =  7'b1100000;     //295pi/512
   m_cos[295]  =  7'b0000011;     //295pi/512
   m_sin[296]  =  7'b1100000;     //296pi/512
   m_cos[296]  =  7'b0000011;     //296pi/512
   m_sin[297]  =  7'b1100000;     //297pi/512
   m_cos[297]  =  7'b0000011;     //297pi/512
   m_sin[298]  =  7'b1100000;     //298pi/512
   m_cos[298]  =  7'b0000011;     //298pi/512
   m_sin[299]  =  7'b1100000;     //299pi/512
   m_cos[299]  =  7'b0000011;     //299pi/512
   m_sin[300]  =  7'b1100000;     //300pi/512
   m_cos[300]  =  7'b0000011;     //300pi/512
   m_sin[301]  =  7'b1100000;     //301pi/512
   m_cos[301]  =  7'b0000010;     //301pi/512
   m_sin[302]  =  7'b1100000;     //302pi/512
   m_cos[302]  =  7'b0000010;     //302pi/512
   m_sin[303]  =  7'b1100000;     //303pi/512
   m_cos[303]  =  7'b0000010;     //303pi/512
   m_sin[304]  =  7'b1100000;     //304pi/512
   m_cos[304]  =  7'b0000010;     //304pi/512
   m_sin[305]  =  7'b1100000;     //305pi/512
   m_cos[305]  =  7'b0000010;     //305pi/512
   m_sin[306]  =  7'b1100000;     //306pi/512
   m_cos[306]  =  7'b0000010;     //306pi/512
   m_sin[307]  =  7'b1100000;     //307pi/512
   m_cos[307]  =  7'b0000010;     //307pi/512
   m_sin[308]  =  7'b1100000;     //308pi/512
   m_cos[308]  =  7'b0000001;     //308pi/512
   m_sin[309]  =  7'b1100000;     //309pi/512
   m_cos[309]  =  7'b0000001;     //309pi/512
   m_sin[310]  =  7'b1100000;     //310pi/512
   m_cos[310]  =  7'b0000001;     //310pi/512
   m_sin[311]  =  7'b1100000;     //311pi/512
   m_cos[311]  =  7'b0000001;     //311pi/512
   m_sin[312]  =  7'b1100000;     //312pi/512
   m_cos[312]  =  7'b0000001;     //312pi/512
   m_sin[313]  =  7'b1100000;     //313pi/512
   m_cos[313]  =  7'b0000001;     //313pi/512
   m_sin[314]  =  7'b1100000;     //314pi/512
   m_cos[314]  =  7'b0000000;     //314pi/512
   m_sin[315]  =  7'b1100000;     //315pi/512
   m_cos[315]  =  7'b0000000;     //315pi/512
   m_sin[316]  =  7'b1100000;     //316pi/512
   m_cos[316]  =  7'b0000000;     //316pi/512
   m_sin[317]  =  7'b1100000;     //317pi/512
   m_cos[317]  =  7'b0000000;     //317pi/512
   m_sin[318]  =  7'b1100000;     //318pi/512
   m_cos[318]  =  7'b0000000;     //318pi/512
   m_sin[319]  =  7'b1100000;     //319pi/512
   m_cos[319]  =  7'b0000000;     //319pi/512
   m_sin[320]  =  7'b1100000;     //320pi/512
   m_cos[320]  =  7'b0000000;     //320pi/512
   m_sin[321]  =  7'b1100000;     //321pi/512
   m_cos[321]  =  7'b0000000;     //321pi/512
   m_sin[322]  =  7'b1100000;     //322pi/512
   m_cos[322]  =  7'b0000000;     //322pi/512
   m_sin[323]  =  7'b1100000;     //323pi/512
   m_cos[323]  =  7'b0000000;     //323pi/512
   m_sin[324]  =  7'b1100000;     //324pi/512
   m_cos[324]  =  7'b1111111;     //324pi/512
   m_sin[325]  =  7'b1100000;     //325pi/512
   m_cos[325]  =  7'b1111111;     //325pi/512
   m_sin[326]  =  7'b1100000;     //326pi/512
   m_cos[326]  =  7'b1111111;     //326pi/512
   m_sin[327]  =  7'b1100000;     //327pi/512
   m_cos[327]  =  7'b1111111;     //327pi/512
   m_sin[328]  =  7'b1100000;     //328pi/512
   m_cos[328]  =  7'b1111111;     //328pi/512
   m_sin[329]  =  7'b1100000;     //329pi/512
   m_cos[329]  =  7'b1111111;     //329pi/512
   m_sin[330]  =  7'b1100000;     //330pi/512
   m_cos[330]  =  7'b1111110;     //330pi/512
   m_sin[331]  =  7'b1100000;     //331pi/512
   m_cos[331]  =  7'b1111110;     //331pi/512
   m_sin[332]  =  7'b1100000;     //332pi/512
   m_cos[332]  =  7'b1111110;     //332pi/512
   m_sin[333]  =  7'b1100000;     //333pi/512
   m_cos[333]  =  7'b1111110;     //333pi/512
   m_sin[334]  =  7'b1100000;     //334pi/512
   m_cos[334]  =  7'b1111110;     //334pi/512
   m_sin[335]  =  7'b1100000;     //335pi/512
   m_cos[335]  =  7'b1111110;     //335pi/512
   m_sin[336]  =  7'b1100000;     //336pi/512
   m_cos[336]  =  7'b1111101;     //336pi/512
   m_sin[337]  =  7'b1100000;     //337pi/512
   m_cos[337]  =  7'b1111101;     //337pi/512
   m_sin[338]  =  7'b1100000;     //338pi/512
   m_cos[338]  =  7'b1111101;     //338pi/512
   m_sin[339]  =  7'b1100000;     //339pi/512
   m_cos[339]  =  7'b1111101;     //339pi/512
   m_sin[340]  =  7'b1100000;     //340pi/512
   m_cos[340]  =  7'b1111101;     //340pi/512
   m_sin[341]  =  7'b1100000;     //341pi/512
   m_cos[341]  =  7'b1111101;     //341pi/512
   m_sin[342]  =  7'b1100000;     //342pi/512
   m_cos[342]  =  7'b1111101;     //342pi/512
   m_sin[343]  =  7'b1100000;     //343pi/512
   m_cos[343]  =  7'b1111100;     //343pi/512
   m_sin[344]  =  7'b1100000;     //344pi/512
   m_cos[344]  =  7'b1111100;     //344pi/512
   m_sin[345]  =  7'b1100000;     //345pi/512
   m_cos[345]  =  7'b1111100;     //345pi/512
   m_sin[346]  =  7'b1100000;     //346pi/512
   m_cos[346]  =  7'b1111100;     //346pi/512
   m_sin[347]  =  7'b1100000;     //347pi/512
   m_cos[347]  =  7'b1111100;     //347pi/512
   m_sin[348]  =  7'b1100000;     //348pi/512
   m_cos[348]  =  7'b1111100;     //348pi/512
   m_sin[349]  =  7'b1100000;     //349pi/512
   m_cos[349]  =  7'b1111011;     //349pi/512
   m_sin[350]  =  7'b1100000;     //350pi/512
   m_cos[350]  =  7'b1111011;     //350pi/512
   m_sin[351]  =  7'b1100000;     //351pi/512
   m_cos[351]  =  7'b1111011;     //351pi/512
   m_sin[352]  =  7'b1100000;     //352pi/512
   m_cos[352]  =  7'b1111011;     //352pi/512
   m_sin[353]  =  7'b1100000;     //353pi/512
   m_cos[353]  =  7'b1111011;     //353pi/512
   m_sin[354]  =  7'b1100000;     //354pi/512
   m_cos[354]  =  7'b1111011;     //354pi/512
   m_sin[355]  =  7'b1100000;     //355pi/512
   m_cos[355]  =  7'b1111011;     //355pi/512
   m_sin[356]  =  7'b1100000;     //356pi/512
   m_cos[356]  =  7'b1111010;     //356pi/512
   m_sin[357]  =  7'b1100001;     //357pi/512
   m_cos[357]  =  7'b1111010;     //357pi/512
   m_sin[358]  =  7'b1100001;     //358pi/512
   m_cos[358]  =  7'b1111010;     //358pi/512
   m_sin[359]  =  7'b1100001;     //359pi/512
   m_cos[359]  =  7'b1111010;     //359pi/512
   m_sin[360]  =  7'b1100001;     //360pi/512
   m_cos[360]  =  7'b1111010;     //360pi/512
   m_sin[361]  =  7'b1100001;     //361pi/512
   m_cos[361]  =  7'b1111010;     //361pi/512
   m_sin[362]  =  7'b1100001;     //362pi/512
   m_cos[362]  =  7'b1111001;     //362pi/512
   m_sin[363]  =  7'b1100001;     //363pi/512
   m_cos[363]  =  7'b1111001;     //363pi/512
   m_sin[364]  =  7'b1100001;     //364pi/512
   m_cos[364]  =  7'b1111001;     //364pi/512
   m_sin[365]  =  7'b1100001;     //365pi/512
   m_cos[365]  =  7'b1111001;     //365pi/512
   m_sin[366]  =  7'b1100001;     //366pi/512
   m_cos[366]  =  7'b1111001;     //366pi/512
   m_sin[367]  =  7'b1100001;     //367pi/512
   m_cos[367]  =  7'b1111001;     //367pi/512
   m_sin[368]  =  7'b1100001;     //368pi/512
   m_cos[368]  =  7'b1111001;     //368pi/512
   m_sin[369]  =  7'b1100001;     //369pi/512
   m_cos[369]  =  7'b1111000;     //369pi/512
   m_sin[370]  =  7'b1100001;     //370pi/512
   m_cos[370]  =  7'b1111000;     //370pi/512
   m_sin[371]  =  7'b1100001;     //371pi/512
   m_cos[371]  =  7'b1111000;     //371pi/512
   m_sin[372]  =  7'b1100001;     //372pi/512
   m_cos[372]  =  7'b1111000;     //372pi/512
   m_sin[373]  =  7'b1100001;     //373pi/512
   m_cos[373]  =  7'b1111000;     //373pi/512
   m_sin[374]  =  7'b1100001;     //374pi/512
   m_cos[374]  =  7'b1111000;     //374pi/512
   m_sin[375]  =  7'b1100001;     //375pi/512
   m_cos[375]  =  7'b1110111;     //375pi/512
   m_sin[376]  =  7'b1100001;     //376pi/512
   m_cos[376]  =  7'b1110111;     //376pi/512
   m_sin[377]  =  7'b1100001;     //377pi/512
   m_cos[377]  =  7'b1110111;     //377pi/512
   m_sin[378]  =  7'b1100001;     //378pi/512
   m_cos[378]  =  7'b1110111;     //378pi/512
   m_sin[379]  =  7'b1100001;     //379pi/512
   m_cos[379]  =  7'b1110111;     //379pi/512
   m_sin[380]  =  7'b1100001;     //380pi/512
   m_cos[380]  =  7'b1110111;     //380pi/512
   m_sin[381]  =  7'b1100001;     //381pi/512
   m_cos[381]  =  7'b1110111;     //381pi/512
   m_sin[382]  =  7'b1100001;     //382pi/512
   m_cos[382]  =  7'b1110110;     //382pi/512
   m_sin[383]  =  7'b1100010;     //383pi/512
   m_cos[383]  =  7'b1110110;     //383pi/512
   m_sin[384]  =  7'b1100010;     //384pi/512
   m_cos[384]  =  7'b1110110;     //384pi/512
   m_sin[385]  =  7'b1100010;     //385pi/512
   m_cos[385]  =  7'b1110110;     //385pi/512
   m_sin[386]  =  7'b1100010;     //386pi/512
   m_cos[386]  =  7'b1110110;     //386pi/512
   m_sin[387]  =  7'b1100010;     //387pi/512
   m_cos[387]  =  7'b1110110;     //387pi/512
   m_sin[388]  =  7'b1100010;     //388pi/512
   m_cos[388]  =  7'b1110110;     //388pi/512
   m_sin[389]  =  7'b1100010;     //389pi/512
   m_cos[389]  =  7'b1110101;     //389pi/512
   m_sin[390]  =  7'b1100010;     //390pi/512
   m_cos[390]  =  7'b1110101;     //390pi/512
   m_sin[391]  =  7'b1100010;     //391pi/512
   m_cos[391]  =  7'b1110101;     //391pi/512
   m_sin[392]  =  7'b1100010;     //392pi/512
   m_cos[392]  =  7'b1110101;     //392pi/512
   m_sin[393]  =  7'b1100010;     //393pi/512
   m_cos[393]  =  7'b1110101;     //393pi/512
   m_sin[394]  =  7'b1100010;     //394pi/512
   m_cos[394]  =  7'b1110101;     //394pi/512
   m_sin[395]  =  7'b1100010;     //395pi/512
   m_cos[395]  =  7'b1110100;     //395pi/512
   m_sin[396]  =  7'b1100010;     //396pi/512
   m_cos[396]  =  7'b1110100;     //396pi/512
   m_sin[397]  =  7'b1100010;     //397pi/512
   m_cos[397]  =  7'b1110100;     //397pi/512
   m_sin[398]  =  7'b1100010;     //398pi/512
   m_cos[398]  =  7'b1110100;     //398pi/512
   m_sin[399]  =  7'b1100010;     //399pi/512
   m_cos[399]  =  7'b1110100;     //399pi/512
   m_sin[400]  =  7'b1100010;     //400pi/512
   m_cos[400]  =  7'b1110100;     //400pi/512
   m_sin[401]  =  7'b1100010;     //401pi/512
   m_cos[401]  =  7'b1110100;     //401pi/512
   m_sin[402]  =  7'b1100011;     //402pi/512
   m_cos[402]  =  7'b1110011;     //402pi/512
   m_sin[403]  =  7'b1100011;     //403pi/512
   m_cos[403]  =  7'b1110011;     //403pi/512
   m_sin[404]  =  7'b1100011;     //404pi/512
   m_cos[404]  =  7'b1110011;     //404pi/512
   m_sin[405]  =  7'b1100011;     //405pi/512
   m_cos[405]  =  7'b1110011;     //405pi/512
   m_sin[406]  =  7'b1100011;     //406pi/512
   m_cos[406]  =  7'b1110011;     //406pi/512
   m_sin[407]  =  7'b1100011;     //407pi/512
   m_cos[407]  =  7'b1110011;     //407pi/512
   m_sin[408]  =  7'b1100011;     //408pi/512
   m_cos[408]  =  7'b1110011;     //408pi/512
   m_sin[409]  =  7'b1100011;     //409pi/512
   m_cos[409]  =  7'b1110010;     //409pi/512
   m_sin[410]  =  7'b1100011;     //410pi/512
   m_cos[410]  =  7'b1110010;     //410pi/512
   m_sin[411]  =  7'b1100011;     //411pi/512
   m_cos[411]  =  7'b1110010;     //411pi/512
   m_sin[412]  =  7'b1100011;     //412pi/512
   m_cos[412]  =  7'b1110010;     //412pi/512
   m_sin[413]  =  7'b1100011;     //413pi/512
   m_cos[413]  =  7'b1110010;     //413pi/512
   m_sin[414]  =  7'b1100011;     //414pi/512
   m_cos[414]  =  7'b1110010;     //414pi/512
   m_sin[415]  =  7'b1100011;     //415pi/512
   m_cos[415]  =  7'b1110010;     //415pi/512
   m_sin[416]  =  7'b1100011;     //416pi/512
   m_cos[416]  =  7'b1110001;     //416pi/512
   m_sin[417]  =  7'b1100100;     //417pi/512
   m_cos[417]  =  7'b1110001;     //417pi/512
   m_sin[418]  =  7'b1100100;     //418pi/512
   m_cos[418]  =  7'b1110001;     //418pi/512
   m_sin[419]  =  7'b1100100;     //419pi/512
   m_cos[419]  =  7'b1110001;     //419pi/512
   m_sin[420]  =  7'b1100100;     //420pi/512
   m_cos[420]  =  7'b1110001;     //420pi/512
   m_sin[421]  =  7'b1100100;     //421pi/512
   m_cos[421]  =  7'b1110001;     //421pi/512
   m_sin[422]  =  7'b1100100;     //422pi/512
   m_cos[422]  =  7'b1110001;     //422pi/512
   m_sin[423]  =  7'b1100100;     //423pi/512
   m_cos[423]  =  7'b1110001;     //423pi/512
   m_sin[424]  =  7'b1100100;     //424pi/512
   m_cos[424]  =  7'b1110000;     //424pi/512
   m_sin[425]  =  7'b1100100;     //425pi/512
   m_cos[425]  =  7'b1110000;     //425pi/512
   m_sin[426]  =  7'b1100100;     //426pi/512
   m_cos[426]  =  7'b1110000;     //426pi/512
   m_sin[427]  =  7'b1100100;     //427pi/512
   m_cos[427]  =  7'b1110000;     //427pi/512
   m_sin[428]  =  7'b1100100;     //428pi/512
   m_cos[428]  =  7'b1110000;     //428pi/512
   m_sin[429]  =  7'b1100100;     //429pi/512
   m_cos[429]  =  7'b1110000;     //429pi/512
   m_sin[430]  =  7'b1100101;     //430pi/512
   m_cos[430]  =  7'b1110000;     //430pi/512
   m_sin[431]  =  7'b1100101;     //431pi/512
   m_cos[431]  =  7'b1101111;     //431pi/512
   m_sin[432]  =  7'b1100101;     //432pi/512
   m_cos[432]  =  7'b1101111;     //432pi/512
   m_sin[433]  =  7'b1100101;     //433pi/512
   m_cos[433]  =  7'b1101111;     //433pi/512
   m_sin[434]  =  7'b1100101;     //434pi/512
   m_cos[434]  =  7'b1101111;     //434pi/512
   m_sin[435]  =  7'b1100101;     //435pi/512
   m_cos[435]  =  7'b1101111;     //435pi/512
   m_sin[436]  =  7'b1100101;     //436pi/512
   m_cos[436]  =  7'b1101111;     //436pi/512
   m_sin[437]  =  7'b1100101;     //437pi/512
   m_cos[437]  =  7'b1101111;     //437pi/512
   m_sin[438]  =  7'b1100101;     //438pi/512
   m_cos[438]  =  7'b1101110;     //438pi/512
   m_sin[439]  =  7'b1100101;     //439pi/512
   m_cos[439]  =  7'b1101110;     //439pi/512
   m_sin[440]  =  7'b1100101;     //440pi/512
   m_cos[440]  =  7'b1101110;     //440pi/512
   m_sin[441]  =  7'b1100101;     //441pi/512
   m_cos[441]  =  7'b1101110;     //441pi/512
   m_sin[442]  =  7'b1100110;     //442pi/512
   m_cos[442]  =  7'b1101110;     //442pi/512
   m_sin[443]  =  7'b1100110;     //443pi/512
   m_cos[443]  =  7'b1101110;     //443pi/512
   m_sin[444]  =  7'b1100110;     //444pi/512
   m_cos[444]  =  7'b1101110;     //444pi/512
   m_sin[445]  =  7'b1100110;     //445pi/512
   m_cos[445]  =  7'b1101110;     //445pi/512
   m_sin[446]  =  7'b1100110;     //446pi/512
   m_cos[446]  =  7'b1101101;     //446pi/512
   m_sin[447]  =  7'b1100110;     //447pi/512
   m_cos[447]  =  7'b1101101;     //447pi/512
   m_sin[448]  =  7'b1100110;     //448pi/512
   m_cos[448]  =  7'b1101101;     //448pi/512
   m_sin[449]  =  7'b1100110;     //449pi/512
   m_cos[449]  =  7'b1101101;     //449pi/512
   m_sin[450]  =  7'b1100110;     //450pi/512
   m_cos[450]  =  7'b1101101;     //450pi/512
   m_sin[451]  =  7'b1100110;     //451pi/512
   m_cos[451]  =  7'b1101101;     //451pi/512
   m_sin[452]  =  7'b1100110;     //452pi/512
   m_cos[452]  =  7'b1101101;     //452pi/512
   m_sin[453]  =  7'b1100111;     //453pi/512
   m_cos[453]  =  7'b1101101;     //453pi/512
   m_sin[454]  =  7'b1100111;     //454pi/512
   m_cos[454]  =  7'b1101100;     //454pi/512
   m_sin[455]  =  7'b1100111;     //455pi/512
   m_cos[455]  =  7'b1101100;     //455pi/512
   m_sin[456]  =  7'b1100111;     //456pi/512
   m_cos[456]  =  7'b1101100;     //456pi/512
   m_sin[457]  =  7'b1100111;     //457pi/512
   m_cos[457]  =  7'b1101100;     //457pi/512
   m_sin[458]  =  7'b1100111;     //458pi/512
   m_cos[458]  =  7'b1101100;     //458pi/512
   m_sin[459]  =  7'b1100111;     //459pi/512
   m_cos[459]  =  7'b1101100;     //459pi/512
   m_sin[460]  =  7'b1100111;     //460pi/512
   m_cos[460]  =  7'b1101100;     //460pi/512
   m_sin[461]  =  7'b1100111;     //461pi/512
   m_cos[461]  =  7'b1101100;     //461pi/512
   m_sin[462]  =  7'b1100111;     //462pi/512
   m_cos[462]  =  7'b1101011;     //462pi/512
   m_sin[463]  =  7'b1101000;     //463pi/512
   m_cos[463]  =  7'b1101011;     //463pi/512
   m_sin[464]  =  7'b1101000;     //464pi/512
   m_cos[464]  =  7'b1101011;     //464pi/512
   m_sin[465]  =  7'b1101000;     //465pi/512
   m_cos[465]  =  7'b1101011;     //465pi/512
   m_sin[466]  =  7'b1101000;     //466pi/512
   m_cos[466]  =  7'b1101011;     //466pi/512
   m_sin[467]  =  7'b1101000;     //467pi/512
   m_cos[467]  =  7'b1101011;     //467pi/512
   m_sin[468]  =  7'b1101000;     //468pi/512
   m_cos[468]  =  7'b1101011;     //468pi/512
   m_sin[469]  =  7'b1101000;     //469pi/512
   m_cos[469]  =  7'b1101011;     //469pi/512
   m_sin[470]  =  7'b1101000;     //470pi/512
   m_cos[470]  =  7'b1101011;     //470pi/512
   m_sin[471]  =  7'b1101000;     //471pi/512
   m_cos[471]  =  7'b1101010;     //471pi/512
   m_sin[472]  =  7'b1101001;     //472pi/512
   m_cos[472]  =  7'b1101010;     //472pi/512
   m_sin[473]  =  7'b1101001;     //473pi/512
   m_cos[473]  =  7'b1101010;     //473pi/512
   m_sin[474]  =  7'b1101001;     //474pi/512
   m_cos[474]  =  7'b1101010;     //474pi/512
   m_sin[475]  =  7'b1101001;     //475pi/512
   m_cos[475]  =  7'b1101010;     //475pi/512
   m_sin[476]  =  7'b1101001;     //476pi/512
   m_cos[476]  =  7'b1101010;     //476pi/512
   m_sin[477]  =  7'b1101001;     //477pi/512
   m_cos[477]  =  7'b1101010;     //477pi/512
   m_sin[478]  =  7'b1101001;     //478pi/512
   m_cos[478]  =  7'b1101010;     //478pi/512
   m_sin[479]  =  7'b1101001;     //479pi/512
   m_cos[479]  =  7'b1101001;     //479pi/512
   m_sin[480]  =  7'b1101001;     //480pi/512
   m_cos[480]  =  7'b1101001;     //480pi/512
   m_sin[481]  =  7'b1101001;     //481pi/512
   m_cos[481]  =  7'b1101001;     //481pi/512
   m_sin[482]  =  7'b1101010;     //482pi/512
   m_cos[482]  =  7'b1101001;     //482pi/512
   m_sin[483]  =  7'b1101010;     //483pi/512
   m_cos[483]  =  7'b1101001;     //483pi/512
   m_sin[484]  =  7'b1101010;     //484pi/512
   m_cos[484]  =  7'b1101001;     //484pi/512
   m_sin[485]  =  7'b1101010;     //485pi/512
   m_cos[485]  =  7'b1101001;     //485pi/512
   m_sin[486]  =  7'b1101010;     //486pi/512
   m_cos[486]  =  7'b1101001;     //486pi/512
   m_sin[487]  =  7'b1101010;     //487pi/512
   m_cos[487]  =  7'b1101001;     //487pi/512
   m_sin[488]  =  7'b1101010;     //488pi/512
   m_cos[488]  =  7'b1101001;     //488pi/512
   m_sin[489]  =  7'b1101010;     //489pi/512
   m_cos[489]  =  7'b1101000;     //489pi/512
   m_sin[490]  =  7'b1101011;     //490pi/512
   m_cos[490]  =  7'b1101000;     //490pi/512
   m_sin[491]  =  7'b1101011;     //491pi/512
   m_cos[491]  =  7'b1101000;     //491pi/512
   m_sin[492]  =  7'b1101011;     //492pi/512
   m_cos[492]  =  7'b1101000;     //492pi/512
   m_sin[493]  =  7'b1101011;     //493pi/512
   m_cos[493]  =  7'b1101000;     //493pi/512
   m_sin[494]  =  7'b1101011;     //494pi/512
   m_cos[494]  =  7'b1101000;     //494pi/512
   m_sin[495]  =  7'b1101011;     //495pi/512
   m_cos[495]  =  7'b1101000;     //495pi/512
   m_sin[496]  =  7'b1101011;     //496pi/512
   m_cos[496]  =  7'b1101000;     //496pi/512
   m_sin[497]  =  7'b1101011;     //497pi/512
   m_cos[497]  =  7'b1101000;     //497pi/512
   m_sin[498]  =  7'b1101011;     //498pi/512
   m_cos[498]  =  7'b1100111;     //498pi/512
   m_sin[499]  =  7'b1101100;     //499pi/512
   m_cos[499]  =  7'b1100111;     //499pi/512
   m_sin[500]  =  7'b1101100;     //500pi/512
   m_cos[500]  =  7'b1100111;     //500pi/512
   m_sin[501]  =  7'b1101100;     //501pi/512
   m_cos[501]  =  7'b1100111;     //501pi/512
   m_sin[502]  =  7'b1101100;     //502pi/512
   m_cos[502]  =  7'b1100111;     //502pi/512
   m_sin[503]  =  7'b1101100;     //503pi/512
   m_cos[503]  =  7'b1100111;     //503pi/512
   m_sin[504]  =  7'b1101100;     //504pi/512
   m_cos[504]  =  7'b1100111;     //504pi/512
   m_sin[505]  =  7'b1101100;     //505pi/512
   m_cos[505]  =  7'b1100111;     //505pi/512
   m_sin[506]  =  7'b1101100;     //506pi/512
   m_cos[506]  =  7'b1100111;     //506pi/512
   m_sin[507]  =  7'b1101101;     //507pi/512
   m_cos[507]  =  7'b1100111;     //507pi/512
   m_sin[508]  =  7'b1101101;     //508pi/512
   m_cos[508]  =  7'b1100110;     //508pi/512
   m_sin[509]  =  7'b1101101;     //509pi/512
   m_cos[509]  =  7'b1100110;     //509pi/512
   m_sin[510]  =  7'b1101101;     //510pi/512
   m_cos[510]  =  7'b1100110;     //510pi/512
   m_sin[511]  =  7'b1101101;     //511pi/512
   m_cos[511]  =  7'b1100110;     //511pi/512
end
endmodule