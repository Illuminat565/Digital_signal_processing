module  TWIDLE_13_bit  #(parameter SIZE = 10, word_length_tw = 13) (
    input            clk,
    input            en_rd,
    input   [10:0]   rd_ptr_angle,
    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );
reg signed [word_length_tw-1:0]  cos  [511:0];
reg signed [word_length_tw-1:0]  sin  [511:0];
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd) begin
                  cos_data           <= cos   [rd_ptr_angle];
                  sin_data           <= sin   [rd_ptr_angle];
             end 
        end
initial begin
   sin[0]  =  13'b0000000000000;     //0pi/512
   cos[0]  =  13'b0100000000000;     //0pi/512
   sin[1]  =  13'b1111111110011;     //1pi/512
   cos[1]  =  13'b0011111111111;     //1pi/512
   sin[2]  =  13'b1111111100111;     //2pi/512
   cos[2]  =  13'b0011111111111;     //2pi/512
   sin[3]  =  13'b1111111011010;     //3pi/512
   cos[3]  =  13'b0011111111111;     //3pi/512
   sin[4]  =  13'b1111111001110;     //4pi/512
   cos[4]  =  13'b0011111111111;     //4pi/512
   sin[5]  =  13'b1111111000001;     //5pi/512
   cos[5]  =  13'b0011111111111;     //5pi/512
   sin[6]  =  13'b1111110110101;     //6pi/512
   cos[6]  =  13'b0011111111110;     //6pi/512
   sin[7]  =  13'b1111110101000;     //7pi/512
   cos[7]  =  13'b0011111111110;     //7pi/512
   sin[8]  =  13'b1111110011100;     //8pi/512
   cos[8]  =  13'b0011111111101;     //8pi/512
   sin[9]  =  13'b1111110001111;     //9pi/512
   cos[9]  =  13'b0011111111100;     //9pi/512
   sin[10]  =  13'b1111110000010;     //10pi/512
   cos[10]  =  13'b0011111111100;     //10pi/512
   sin[11]  =  13'b1111101110110;     //11pi/512
   cos[11]  =  13'b0011111111011;     //11pi/512
   sin[12]  =  13'b1111101101001;     //12pi/512
   cos[12]  =  13'b0011111111010;     //12pi/512
   sin[13]  =  13'b1111101011101;     //13pi/512
   cos[13]  =  13'b0011111111001;     //13pi/512
   sin[14]  =  13'b1111101010000;     //14pi/512
   cos[14]  =  13'b0011111111000;     //14pi/512
   sin[15]  =  13'b1111101000100;     //15pi/512
   cos[15]  =  13'b0011111110111;     //15pi/512
   sin[16]  =  13'b1111100110111;     //16pi/512
   cos[16]  =  13'b0011111110110;     //16pi/512
   sin[17]  =  13'b1111100101011;     //17pi/512
   cos[17]  =  13'b0011111110100;     //17pi/512
   sin[18]  =  13'b1111100011110;     //18pi/512
   cos[18]  =  13'b0011111110011;     //18pi/512
   sin[19]  =  13'b1111100010010;     //19pi/512
   cos[19]  =  13'b0011111110010;     //19pi/512
   sin[20]  =  13'b1111100000101;     //20pi/512
   cos[20]  =  13'b0011111110000;     //20pi/512
   sin[21]  =  13'b1111011111001;     //21pi/512
   cos[21]  =  13'b0011111101111;     //21pi/512
   sin[22]  =  13'b1111011101100;     //22pi/512
   cos[22]  =  13'b0011111101101;     //22pi/512
   sin[23]  =  13'b1111011100000;     //23pi/512
   cos[23]  =  13'b0011111101011;     //23pi/512
   sin[24]  =  13'b1111011010011;     //24pi/512
   cos[24]  =  13'b0011111101001;     //24pi/512
   sin[25]  =  13'b1111011000111;     //25pi/512
   cos[25]  =  13'b0011111100111;     //25pi/512
   sin[26]  =  13'b1111010111011;     //26pi/512
   cos[26]  =  13'b0011111100101;     //26pi/512
   sin[27]  =  13'b1111010101110;     //27pi/512
   cos[27]  =  13'b0011111100011;     //27pi/512
   sin[28]  =  13'b1111010100010;     //28pi/512
   cos[28]  =  13'b0011111100001;     //28pi/512
   sin[29]  =  13'b1111010010101;     //29pi/512
   cos[29]  =  13'b0011111011111;     //29pi/512
   sin[30]  =  13'b1111010001001;     //30pi/512
   cos[30]  =  13'b0011111011101;     //30pi/512
   sin[31]  =  13'b1111001111101;     //31pi/512
   cos[31]  =  13'b0011111011011;     //31pi/512
   sin[32]  =  13'b1111001110000;     //32pi/512
   cos[32]  =  13'b0011111011000;     //32pi/512
   sin[33]  =  13'b1111001100100;     //33pi/512
   cos[33]  =  13'b0011111010110;     //33pi/512
   sin[34]  =  13'b1111001011000;     //34pi/512
   cos[34]  =  13'b0011111010011;     //34pi/512
   sin[35]  =  13'b1111001001100;     //35pi/512
   cos[35]  =  13'b0011111010000;     //35pi/512
   sin[36]  =  13'b1111000111111;     //36pi/512
   cos[36]  =  13'b0011111001110;     //36pi/512
   sin[37]  =  13'b1111000110011;     //37pi/512
   cos[37]  =  13'b0011111001011;     //37pi/512
   sin[38]  =  13'b1111000100111;     //38pi/512
   cos[38]  =  13'b0011111001000;     //38pi/512
   sin[39]  =  13'b1111000011011;     //39pi/512
   cos[39]  =  13'b0011111000101;     //39pi/512
   sin[40]  =  13'b1111000001110;     //40pi/512
   cos[40]  =  13'b0011111000010;     //40pi/512
   sin[41]  =  13'b1111000000010;     //41pi/512
   cos[41]  =  13'b0011110111111;     //41pi/512
   sin[42]  =  13'b1110111110110;     //42pi/512
   cos[42]  =  13'b0011110111100;     //42pi/512
   sin[43]  =  13'b1110111101010;     //43pi/512
   cos[43]  =  13'b0011110111001;     //43pi/512
   sin[44]  =  13'b1110111011110;     //44pi/512
   cos[44]  =  13'b0011110110101;     //44pi/512
   sin[45]  =  13'b1110111010010;     //45pi/512
   cos[45]  =  13'b0011110110010;     //45pi/512
   sin[46]  =  13'b1110111000110;     //46pi/512
   cos[46]  =  13'b0011110101110;     //46pi/512
   sin[47]  =  13'b1110110111010;     //47pi/512
   cos[47]  =  13'b0011110101011;     //47pi/512
   sin[48]  =  13'b1110110101101;     //48pi/512
   cos[48]  =  13'b0011110100111;     //48pi/512
   sin[49]  =  13'b1110110100001;     //49pi/512
   cos[49]  =  13'b0011110100100;     //49pi/512
   sin[50]  =  13'b1110110010101;     //50pi/512
   cos[50]  =  13'b0011110100000;     //50pi/512
   sin[51]  =  13'b1110110001010;     //51pi/512
   cos[51]  =  13'b0011110011100;     //51pi/512
   sin[52]  =  13'b1110101111110;     //52pi/512
   cos[52]  =  13'b0011110011000;     //52pi/512
   sin[53]  =  13'b1110101110010;     //53pi/512
   cos[53]  =  13'b0011110010100;     //53pi/512
   sin[54]  =  13'b1110101100110;     //54pi/512
   cos[54]  =  13'b0011110010000;     //54pi/512
   sin[55]  =  13'b1110101011010;     //55pi/512
   cos[55]  =  13'b0011110001100;     //55pi/512
   sin[56]  =  13'b1110101001110;     //56pi/512
   cos[56]  =  13'b0011110001000;     //56pi/512
   sin[57]  =  13'b1110101000010;     //57pi/512
   cos[57]  =  13'b0011110000100;     //57pi/512
   sin[58]  =  13'b1110100110110;     //58pi/512
   cos[58]  =  13'b0011101111111;     //58pi/512
   sin[59]  =  13'b1110100101011;     //59pi/512
   cos[59]  =  13'b0011101111011;     //59pi/512
   sin[60]  =  13'b1110100011111;     //60pi/512
   cos[60]  =  13'b0011101110110;     //60pi/512
   sin[61]  =  13'b1110100010011;     //61pi/512
   cos[61]  =  13'b0011101110010;     //61pi/512
   sin[62]  =  13'b1110100001000;     //62pi/512
   cos[62]  =  13'b0011101101101;     //62pi/512
   sin[63]  =  13'b1110011111100;     //63pi/512
   cos[63]  =  13'b0011101101000;     //63pi/512
   sin[64]  =  13'b1110011110000;     //64pi/512
   cos[64]  =  13'b0011101100100;     //64pi/512
   sin[65]  =  13'b1110011100101;     //65pi/512
   cos[65]  =  13'b0011101011111;     //65pi/512
   sin[66]  =  13'b1110011011001;     //66pi/512
   cos[66]  =  13'b0011101011010;     //66pi/512
   sin[67]  =  13'b1110011001110;     //67pi/512
   cos[67]  =  13'b0011101010101;     //67pi/512
   sin[68]  =  13'b1110011000010;     //68pi/512
   cos[68]  =  13'b0011101010000;     //68pi/512
   sin[69]  =  13'b1110010110111;     //69pi/512
   cos[69]  =  13'b0011101001011;     //69pi/512
   sin[70]  =  13'b1110010101011;     //70pi/512
   cos[70]  =  13'b0011101000101;     //70pi/512
   sin[71]  =  13'b1110010100000;     //71pi/512
   cos[71]  =  13'b0011101000000;     //71pi/512
   sin[72]  =  13'b1110010010100;     //72pi/512
   cos[72]  =  13'b0011100111011;     //72pi/512
   sin[73]  =  13'b1110010001001;     //73pi/512
   cos[73]  =  13'b0011100110101;     //73pi/512
   sin[74]  =  13'b1110001111110;     //74pi/512
   cos[74]  =  13'b0011100110000;     //74pi/512
   sin[75]  =  13'b1110001110010;     //75pi/512
   cos[75]  =  13'b0011100101010;     //75pi/512
   sin[76]  =  13'b1110001100111;     //76pi/512
   cos[76]  =  13'b0011100100101;     //76pi/512
   sin[77]  =  13'b1110001011100;     //77pi/512
   cos[77]  =  13'b0011100011111;     //77pi/512
   sin[78]  =  13'b1110001010001;     //78pi/512
   cos[78]  =  13'b0011100011001;     //78pi/512
   sin[79]  =  13'b1110001000110;     //79pi/512
   cos[79]  =  13'b0011100010100;     //79pi/512
   sin[80]  =  13'b1110000111011;     //80pi/512
   cos[80]  =  13'b0011100001110;     //80pi/512
   sin[81]  =  13'b1110000110000;     //81pi/512
   cos[81]  =  13'b0011100001000;     //81pi/512
   sin[82]  =  13'b1110000100100;     //82pi/512
   cos[82]  =  13'b0011100000010;     //82pi/512
   sin[83]  =  13'b1110000011001;     //83pi/512
   cos[83]  =  13'b0011011111100;     //83pi/512
   sin[84]  =  13'b1110000001111;     //84pi/512
   cos[84]  =  13'b0011011110101;     //84pi/512
   sin[85]  =  13'b1110000000100;     //85pi/512
   cos[85]  =  13'b0011011101111;     //85pi/512
   sin[86]  =  13'b1101111111001;     //86pi/512
   cos[86]  =  13'b0011011101001;     //86pi/512
   sin[87]  =  13'b1101111101110;     //87pi/512
   cos[87]  =  13'b0011011100011;     //87pi/512
   sin[88]  =  13'b1101111100011;     //88pi/512
   cos[88]  =  13'b0011011011100;     //88pi/512
   sin[89]  =  13'b1101111011000;     //89pi/512
   cos[89]  =  13'b0011011010110;     //89pi/512
   sin[90]  =  13'b1101111001110;     //90pi/512
   cos[90]  =  13'b0011011001111;     //90pi/512
   sin[91]  =  13'b1101111000011;     //91pi/512
   cos[91]  =  13'b0011011001000;     //91pi/512
   sin[92]  =  13'b1101110111000;     //92pi/512
   cos[92]  =  13'b0011011000010;     //92pi/512
   sin[93]  =  13'b1101110101110;     //93pi/512
   cos[93]  =  13'b0011010111011;     //93pi/512
   sin[94]  =  13'b1101110100011;     //94pi/512
   cos[94]  =  13'b0011010110100;     //94pi/512
   sin[95]  =  13'b1101110011001;     //95pi/512
   cos[95]  =  13'b0011010101101;     //95pi/512
   sin[96]  =  13'b1101110001110;     //96pi/512
   cos[96]  =  13'b0011010100110;     //96pi/512
   sin[97]  =  13'b1101110000100;     //97pi/512
   cos[97]  =  13'b0011010011111;     //97pi/512
   sin[98]  =  13'b1101101111001;     //98pi/512
   cos[98]  =  13'b0011010011000;     //98pi/512
   sin[99]  =  13'b1101101101111;     //99pi/512
   cos[99]  =  13'b0011010010001;     //99pi/512
   sin[100]  =  13'b1101101100101;     //100pi/512
   cos[100]  =  13'b0011010001010;     //100pi/512
   sin[101]  =  13'b1101101011010;     //101pi/512
   cos[101]  =  13'b0011010000011;     //101pi/512
   sin[102]  =  13'b1101101010000;     //102pi/512
   cos[102]  =  13'b0011001111011;     //102pi/512
   sin[103]  =  13'b1101101000110;     //103pi/512
   cos[103]  =  13'b0011001110100;     //103pi/512
   sin[104]  =  13'b1101100111100;     //104pi/512
   cos[104]  =  13'b0011001101100;     //104pi/512
   sin[105]  =  13'b1101100110010;     //105pi/512
   cos[105]  =  13'b0011001100101;     //105pi/512
   sin[106]  =  13'b1101100101000;     //106pi/512
   cos[106]  =  13'b0011001011101;     //106pi/512
   sin[107]  =  13'b1101100011110;     //107pi/512
   cos[107]  =  13'b0011001010110;     //107pi/512
   sin[108]  =  13'b1101100010100;     //108pi/512
   cos[108]  =  13'b0011001001110;     //108pi/512
   sin[109]  =  13'b1101100001010;     //109pi/512
   cos[109]  =  13'b0011001000110;     //109pi/512
   sin[110]  =  13'b1101100000000;     //110pi/512
   cos[110]  =  13'b0011000111110;     //110pi/512
   sin[111]  =  13'b1101011110111;     //111pi/512
   cos[111]  =  13'b0011000110111;     //111pi/512
   sin[112]  =  13'b1101011101101;     //112pi/512
   cos[112]  =  13'b0011000101111;     //112pi/512
   sin[113]  =  13'b1101011100011;     //113pi/512
   cos[113]  =  13'b0011000100111;     //113pi/512
   sin[114]  =  13'b1101011011001;     //114pi/512
   cos[114]  =  13'b0011000011111;     //114pi/512
   sin[115]  =  13'b1101011010000;     //115pi/512
   cos[115]  =  13'b0011000010110;     //115pi/512
   sin[116]  =  13'b1101011000110;     //116pi/512
   cos[116]  =  13'b0011000001110;     //116pi/512
   sin[117]  =  13'b1101010111101;     //117pi/512
   cos[117]  =  13'b0011000000110;     //117pi/512
   sin[118]  =  13'b1101010110011;     //118pi/512
   cos[118]  =  13'b0010111111110;     //118pi/512
   sin[119]  =  13'b1101010101010;     //119pi/512
   cos[119]  =  13'b0010111110101;     //119pi/512
   sin[120]  =  13'b1101010100001;     //120pi/512
   cos[120]  =  13'b0010111101101;     //120pi/512
   sin[121]  =  13'b1101010010111;     //121pi/512
   cos[121]  =  13'b0010111100101;     //121pi/512
   sin[122]  =  13'b1101010001110;     //122pi/512
   cos[122]  =  13'b0010111011100;     //122pi/512
   sin[123]  =  13'b1101010000101;     //123pi/512
   cos[123]  =  13'b0010111010011;     //123pi/512
   sin[124]  =  13'b1101001111100;     //124pi/512
   cos[124]  =  13'b0010111001011;     //124pi/512
   sin[125]  =  13'b1101001110011;     //125pi/512
   cos[125]  =  13'b0010111000010;     //125pi/512
   sin[126]  =  13'b1101001101010;     //126pi/512
   cos[126]  =  13'b0010110111001;     //126pi/512
   sin[127]  =  13'b1101001100001;     //127pi/512
   cos[127]  =  13'b0010110110001;     //127pi/512
   sin[128]  =  13'b1101001011000;     //128pi/512
   cos[128]  =  13'b0010110101000;     //128pi/512
   sin[129]  =  13'b1101001001111;     //129pi/512
   cos[129]  =  13'b0010110011111;     //129pi/512
   sin[130]  =  13'b1101001000110;     //130pi/512
   cos[130]  =  13'b0010110010110;     //130pi/512
   sin[131]  =  13'b1101000111101;     //131pi/512
   cos[131]  =  13'b0010110001101;     //131pi/512
   sin[132]  =  13'b1101000110101;     //132pi/512
   cos[132]  =  13'b0010110000100;     //132pi/512
   sin[133]  =  13'b1101000101100;     //133pi/512
   cos[133]  =  13'b0010101111011;     //133pi/512
   sin[134]  =  13'b1101000100100;     //134pi/512
   cos[134]  =  13'b0010101110001;     //134pi/512
   sin[135]  =  13'b1101000011011;     //135pi/512
   cos[135]  =  13'b0010101101000;     //135pi/512
   sin[136]  =  13'b1101000010011;     //136pi/512
   cos[136]  =  13'b0010101011111;     //136pi/512
   sin[137]  =  13'b1101000001010;     //137pi/512
   cos[137]  =  13'b0010101010110;     //137pi/512
   sin[138]  =  13'b1101000000010;     //138pi/512
   cos[138]  =  13'b0010101001100;     //138pi/512
   sin[139]  =  13'b1100111111001;     //139pi/512
   cos[139]  =  13'b0010101000011;     //139pi/512
   sin[140]  =  13'b1100111110001;     //140pi/512
   cos[140]  =  13'b0010100111001;     //140pi/512
   sin[141]  =  13'b1100111101001;     //141pi/512
   cos[141]  =  13'b0010100110000;     //141pi/512
   sin[142]  =  13'b1100111100001;     //142pi/512
   cos[142]  =  13'b0010100100110;     //142pi/512
   sin[143]  =  13'b1100111011001;     //143pi/512
   cos[143]  =  13'b0010100011100;     //143pi/512
   sin[144]  =  13'b1100111010001;     //144pi/512
   cos[144]  =  13'b0010100010011;     //144pi/512
   sin[145]  =  13'b1100111001001;     //145pi/512
   cos[145]  =  13'b0010100001001;     //145pi/512
   sin[146]  =  13'b1100111000001;     //146pi/512
   cos[146]  =  13'b0010011111111;     //146pi/512
   sin[147]  =  13'b1100110111001;     //147pi/512
   cos[147]  =  13'b0010011110101;     //147pi/512
   sin[148]  =  13'b1100110110001;     //148pi/512
   cos[148]  =  13'b0010011101011;     //148pi/512
   sin[149]  =  13'b1100110101010;     //149pi/512
   cos[149]  =  13'b0010011100010;     //149pi/512
   sin[150]  =  13'b1100110100010;     //150pi/512
   cos[150]  =  13'b0010011011000;     //150pi/512
   sin[151]  =  13'b1100110011011;     //151pi/512
   cos[151]  =  13'b0010011001110;     //151pi/512
   sin[152]  =  13'b1100110010011;     //152pi/512
   cos[152]  =  13'b0010011000011;     //152pi/512
   sin[153]  =  13'b1100110001100;     //153pi/512
   cos[153]  =  13'b0010010111001;     //153pi/512
   sin[154]  =  13'b1100110000100;     //154pi/512
   cos[154]  =  13'b0010010101111;     //154pi/512
   sin[155]  =  13'b1100101111101;     //155pi/512
   cos[155]  =  13'b0010010100101;     //155pi/512
   sin[156]  =  13'b1100101110110;     //156pi/512
   cos[156]  =  13'b0010010011011;     //156pi/512
   sin[157]  =  13'b1100101101110;     //157pi/512
   cos[157]  =  13'b0010010010000;     //157pi/512
   sin[158]  =  13'b1100101100111;     //158pi/512
   cos[158]  =  13'b0010010000110;     //158pi/512
   sin[159]  =  13'b1100101100000;     //159pi/512
   cos[159]  =  13'b0010001111100;     //159pi/512
   sin[160]  =  13'b1100101011001;     //160pi/512
   cos[160]  =  13'b0010001110001;     //160pi/512
   sin[161]  =  13'b1100101010010;     //161pi/512
   cos[161]  =  13'b0010001100111;     //161pi/512
   sin[162]  =  13'b1100101001011;     //162pi/512
   cos[162]  =  13'b0010001011100;     //162pi/512
   sin[163]  =  13'b1100101000100;     //163pi/512
   cos[163]  =  13'b0010001010010;     //163pi/512
   sin[164]  =  13'b1100100111110;     //164pi/512
   cos[164]  =  13'b0010001000111;     //164pi/512
   sin[165]  =  13'b1100100110111;     //165pi/512
   cos[165]  =  13'b0010000111101;     //165pi/512
   sin[166]  =  13'b1100100110000;     //166pi/512
   cos[166]  =  13'b0010000110010;     //166pi/512
   sin[167]  =  13'b1100100101010;     //167pi/512
   cos[167]  =  13'b0010000100111;     //167pi/512
   sin[168]  =  13'b1100100100011;     //168pi/512
   cos[168]  =  13'b0010000011100;     //168pi/512
   sin[169]  =  13'b1100100011101;     //169pi/512
   cos[169]  =  13'b0010000010010;     //169pi/512
   sin[170]  =  13'b1100100010111;     //170pi/512
   cos[170]  =  13'b0010000000111;     //170pi/512
   sin[171]  =  13'b1100100010000;     //171pi/512
   cos[171]  =  13'b0001111111100;     //171pi/512
   sin[172]  =  13'b1100100001010;     //172pi/512
   cos[172]  =  13'b0001111110001;     //172pi/512
   sin[173]  =  13'b1100100000100;     //173pi/512
   cos[173]  =  13'b0001111100110;     //173pi/512
   sin[174]  =  13'b1100011111110;     //174pi/512
   cos[174]  =  13'b0001111011011;     //174pi/512
   sin[175]  =  13'b1100011111000;     //175pi/512
   cos[175]  =  13'b0001111010000;     //175pi/512
   sin[176]  =  13'b1100011110010;     //176pi/512
   cos[176]  =  13'b0001111000101;     //176pi/512
   sin[177]  =  13'b1100011101100;     //177pi/512
   cos[177]  =  13'b0001110111010;     //177pi/512
   sin[178]  =  13'b1100011100110;     //178pi/512
   cos[178]  =  13'b0001110101111;     //178pi/512
   sin[179]  =  13'b1100011100000;     //179pi/512
   cos[179]  =  13'b0001110100100;     //179pi/512
   sin[180]  =  13'b1100011011011;     //180pi/512
   cos[180]  =  13'b0001110011000;     //180pi/512
   sin[181]  =  13'b1100011010101;     //181pi/512
   cos[181]  =  13'b0001110001101;     //181pi/512
   sin[182]  =  13'b1100011010000;     //182pi/512
   cos[182]  =  13'b0001110000010;     //182pi/512
   sin[183]  =  13'b1100011001010;     //183pi/512
   cos[183]  =  13'b0001101110110;     //183pi/512
   sin[184]  =  13'b1100011000101;     //184pi/512
   cos[184]  =  13'b0001101101011;     //184pi/512
   sin[185]  =  13'b1100010111111;     //185pi/512
   cos[185]  =  13'b0001101100000;     //185pi/512
   sin[186]  =  13'b1100010111010;     //186pi/512
   cos[186]  =  13'b0001101010100;     //186pi/512
   sin[187]  =  13'b1100010110101;     //187pi/512
   cos[187]  =  13'b0001101001001;     //187pi/512
   sin[188]  =  13'b1100010110000;     //188pi/512
   cos[188]  =  13'b0001100111101;     //188pi/512
   sin[189]  =  13'b1100010101011;     //189pi/512
   cos[189]  =  13'b0001100110010;     //189pi/512
   sin[190]  =  13'b1100010100110;     //190pi/512
   cos[190]  =  13'b0001100100110;     //190pi/512
   sin[191]  =  13'b1100010100001;     //191pi/512
   cos[191]  =  13'b0001100011011;     //191pi/512
   sin[192]  =  13'b1100010011100;     //192pi/512
   cos[192]  =  13'b0001100001111;     //192pi/512
   sin[193]  =  13'b1100010010111;     //193pi/512
   cos[193]  =  13'b0001100000100;     //193pi/512
   sin[194]  =  13'b1100010010010;     //194pi/512
   cos[194]  =  13'b0001011111000;     //194pi/512
   sin[195]  =  13'b1100010001110;     //195pi/512
   cos[195]  =  13'b0001011101100;     //195pi/512
   sin[196]  =  13'b1100010001001;     //196pi/512
   cos[196]  =  13'b0001011100001;     //196pi/512
   sin[197]  =  13'b1100010000101;     //197pi/512
   cos[197]  =  13'b0001011010101;     //197pi/512
   sin[198]  =  13'b1100010000000;     //198pi/512
   cos[198]  =  13'b0001011001001;     //198pi/512
   sin[199]  =  13'b1100001111100;     //199pi/512
   cos[199]  =  13'b0001010111101;     //199pi/512
   sin[200]  =  13'b1100001111000;     //200pi/512
   cos[200]  =  13'b0001010110001;     //200pi/512
   sin[201]  =  13'b1100001110100;     //201pi/512
   cos[201]  =  13'b0001010100110;     //201pi/512
   sin[202]  =  13'b1100001101111;     //202pi/512
   cos[202]  =  13'b0001010011010;     //202pi/512
   sin[203]  =  13'b1100001101011;     //203pi/512
   cos[203]  =  13'b0001010001110;     //203pi/512
   sin[204]  =  13'b1100001100111;     //204pi/512
   cos[204]  =  13'b0001010000010;     //204pi/512
   sin[205]  =  13'b1100001100011;     //205pi/512
   cos[205]  =  13'b0001001110110;     //205pi/512
   sin[206]  =  13'b1100001100000;     //206pi/512
   cos[206]  =  13'b0001001101010;     //206pi/512
   sin[207]  =  13'b1100001011100;     //207pi/512
   cos[207]  =  13'b0001001011110;     //207pi/512
   sin[208]  =  13'b1100001011000;     //208pi/512
   cos[208]  =  13'b0001001010010;     //208pi/512
   sin[209]  =  13'b1100001010101;     //209pi/512
   cos[209]  =  13'b0001001000110;     //209pi/512
   sin[210]  =  13'b1100001010001;     //210pi/512
   cos[210]  =  13'b0001000111010;     //210pi/512
   sin[211]  =  13'b1100001001110;     //211pi/512
   cos[211]  =  13'b0001000101110;     //211pi/512
   sin[212]  =  13'b1100001001010;     //212pi/512
   cos[212]  =  13'b0001000100010;     //212pi/512
   sin[213]  =  13'b1100001000111;     //213pi/512
   cos[213]  =  13'b0001000010110;     //213pi/512
   sin[214]  =  13'b1100001000100;     //214pi/512
   cos[214]  =  13'b0001000001001;     //214pi/512
   sin[215]  =  13'b1100001000000;     //215pi/512
   cos[215]  =  13'b0000111111101;     //215pi/512
   sin[216]  =  13'b1100000111101;     //216pi/512
   cos[216]  =  13'b0000111110001;     //216pi/512
   sin[217]  =  13'b1100000111010;     //217pi/512
   cos[217]  =  13'b0000111100101;     //217pi/512
   sin[218]  =  13'b1100000110111;     //218pi/512
   cos[218]  =  13'b0000111011001;     //218pi/512
   sin[219]  =  13'b1100000110101;     //219pi/512
   cos[219]  =  13'b0000111001100;     //219pi/512
   sin[220]  =  13'b1100000110010;     //220pi/512
   cos[220]  =  13'b0000111000000;     //220pi/512
   sin[221]  =  13'b1100000101111;     //221pi/512
   cos[221]  =  13'b0000110110100;     //221pi/512
   sin[222]  =  13'b1100000101100;     //222pi/512
   cos[222]  =  13'b0000110101000;     //222pi/512
   sin[223]  =  13'b1100000101010;     //223pi/512
   cos[223]  =  13'b0000110011011;     //223pi/512
   sin[224]  =  13'b1100000100111;     //224pi/512
   cos[224]  =  13'b0000110001111;     //224pi/512
   sin[225]  =  13'b1100000100101;     //225pi/512
   cos[225]  =  13'b0000110000011;     //225pi/512
   sin[226]  =  13'b1100000100011;     //226pi/512
   cos[226]  =  13'b0000101110110;     //226pi/512
   sin[227]  =  13'b1100000100000;     //227pi/512
   cos[227]  =  13'b0000101101010;     //227pi/512
   sin[228]  =  13'b1100000011110;     //228pi/512
   cos[228]  =  13'b0000101011110;     //228pi/512
   sin[229]  =  13'b1100000011100;     //229pi/512
   cos[229]  =  13'b0000101010001;     //229pi/512
   sin[230]  =  13'b1100000011010;     //230pi/512
   cos[230]  =  13'b0000101000101;     //230pi/512
   sin[231]  =  13'b1100000011000;     //231pi/512
   cos[231]  =  13'b0000100111000;     //231pi/512
   sin[232]  =  13'b1100000010110;     //232pi/512
   cos[232]  =  13'b0000100101100;     //232pi/512
   sin[233]  =  13'b1100000010100;     //233pi/512
   cos[233]  =  13'b0000100100000;     //233pi/512
   sin[234]  =  13'b1100000010011;     //234pi/512
   cos[234]  =  13'b0000100010011;     //234pi/512
   sin[235]  =  13'b1100000010001;     //235pi/512
   cos[235]  =  13'b0000100000111;     //235pi/512
   sin[236]  =  13'b1100000001111;     //236pi/512
   cos[236]  =  13'b0000011111010;     //236pi/512
   sin[237]  =  13'b1100000001110;     //237pi/512
   cos[237]  =  13'b0000011101110;     //237pi/512
   sin[238]  =  13'b1100000001100;     //238pi/512
   cos[238]  =  13'b0000011100001;     //238pi/512
   sin[239]  =  13'b1100000001011;     //239pi/512
   cos[239]  =  13'b0000011010101;     //239pi/512
   sin[240]  =  13'b1100000001010;     //240pi/512
   cos[240]  =  13'b0000011001000;     //240pi/512
   sin[241]  =  13'b1100000001001;     //241pi/512
   cos[241]  =  13'b0000010111100;     //241pi/512
   sin[242]  =  13'b1100000001000;     //242pi/512
   cos[242]  =  13'b0000010101111;     //242pi/512
   sin[243]  =  13'b1100000000111;     //243pi/512
   cos[243]  =  13'b0000010100011;     //243pi/512
   sin[244]  =  13'b1100000000110;     //244pi/512
   cos[244]  =  13'b0000010010110;     //244pi/512
   sin[245]  =  13'b1100000000101;     //245pi/512
   cos[245]  =  13'b0000010001010;     //245pi/512
   sin[246]  =  13'b1100000000100;     //246pi/512
   cos[246]  =  13'b0000001111101;     //246pi/512
   sin[247]  =  13'b1100000000011;     //247pi/512
   cos[247]  =  13'b0000001110001;     //247pi/512
   sin[248]  =  13'b1100000000010;     //248pi/512
   cos[248]  =  13'b0000001100100;     //248pi/512
   sin[249]  =  13'b1100000000010;     //249pi/512
   cos[249]  =  13'b0000001010111;     //249pi/512
   sin[250]  =  13'b1100000000001;     //250pi/512
   cos[250]  =  13'b0000001001011;     //250pi/512
   sin[251]  =  13'b1100000000001;     //251pi/512
   cos[251]  =  13'b0000000111110;     //251pi/512
   sin[252]  =  13'b1100000000001;     //252pi/512
   cos[252]  =  13'b0000000110010;     //252pi/512
   sin[253]  =  13'b1100000000000;     //253pi/512
   cos[253]  =  13'b0000000100101;     //253pi/512
   sin[254]  =  13'b1100000000000;     //254pi/512
   cos[254]  =  13'b0000000011001;     //254pi/512
   sin[255]  =  13'b1100000000000;     //255pi/512
   cos[255]  =  13'b0000000001100;     //255pi/512
   sin[256]  =  13'b1100000000000;     //256pi/512
   cos[256]  =  13'b0000000000000;     //256pi/512
   sin[257]  =  13'b1100000000000;     //257pi/512
   cos[257]  =  13'b1111111110011;     //257pi/512
   sin[258]  =  13'b1100000000000;     //258pi/512
   cos[258]  =  13'b1111111100111;     //258pi/512
   sin[259]  =  13'b1100000000000;     //259pi/512
   cos[259]  =  13'b1111111011010;     //259pi/512
   sin[260]  =  13'b1100000000001;     //260pi/512
   cos[260]  =  13'b1111111001110;     //260pi/512
   sin[261]  =  13'b1100000000001;     //261pi/512
   cos[261]  =  13'b1111111000001;     //261pi/512
   sin[262]  =  13'b1100000000001;     //262pi/512
   cos[262]  =  13'b1111110110101;     //262pi/512
   sin[263]  =  13'b1100000000010;     //263pi/512
   cos[263]  =  13'b1111110101000;     //263pi/512
   sin[264]  =  13'b1100000000010;     //264pi/512
   cos[264]  =  13'b1111110011100;     //264pi/512
   sin[265]  =  13'b1100000000011;     //265pi/512
   cos[265]  =  13'b1111110001111;     //265pi/512
   sin[266]  =  13'b1100000000100;     //266pi/512
   cos[266]  =  13'b1111110000010;     //266pi/512
   sin[267]  =  13'b1100000000101;     //267pi/512
   cos[267]  =  13'b1111101110110;     //267pi/512
   sin[268]  =  13'b1100000000110;     //268pi/512
   cos[268]  =  13'b1111101101001;     //268pi/512
   sin[269]  =  13'b1100000000111;     //269pi/512
   cos[269]  =  13'b1111101011101;     //269pi/512
   sin[270]  =  13'b1100000001000;     //270pi/512
   cos[270]  =  13'b1111101010000;     //270pi/512
   sin[271]  =  13'b1100000001001;     //271pi/512
   cos[271]  =  13'b1111101000100;     //271pi/512
   sin[272]  =  13'b1100000001010;     //272pi/512
   cos[272]  =  13'b1111100110111;     //272pi/512
   sin[273]  =  13'b1100000001011;     //273pi/512
   cos[273]  =  13'b1111100101011;     //273pi/512
   sin[274]  =  13'b1100000001100;     //274pi/512
   cos[274]  =  13'b1111100011110;     //274pi/512
   sin[275]  =  13'b1100000001110;     //275pi/512
   cos[275]  =  13'b1111100010010;     //275pi/512
   sin[276]  =  13'b1100000001111;     //276pi/512
   cos[276]  =  13'b1111100000101;     //276pi/512
   sin[277]  =  13'b1100000010001;     //277pi/512
   cos[277]  =  13'b1111011111001;     //277pi/512
   sin[278]  =  13'b1100000010011;     //278pi/512
   cos[278]  =  13'b1111011101100;     //278pi/512
   sin[279]  =  13'b1100000010100;     //279pi/512
   cos[279]  =  13'b1111011100000;     //279pi/512
   sin[280]  =  13'b1100000010110;     //280pi/512
   cos[280]  =  13'b1111011010011;     //280pi/512
   sin[281]  =  13'b1100000011000;     //281pi/512
   cos[281]  =  13'b1111011000111;     //281pi/512
   sin[282]  =  13'b1100000011010;     //282pi/512
   cos[282]  =  13'b1111010111011;     //282pi/512
   sin[283]  =  13'b1100000011100;     //283pi/512
   cos[283]  =  13'b1111010101110;     //283pi/512
   sin[284]  =  13'b1100000011110;     //284pi/512
   cos[284]  =  13'b1111010100010;     //284pi/512
   sin[285]  =  13'b1100000100000;     //285pi/512
   cos[285]  =  13'b1111010010101;     //285pi/512
   sin[286]  =  13'b1100000100011;     //286pi/512
   cos[286]  =  13'b1111010001001;     //286pi/512
   sin[287]  =  13'b1100000100101;     //287pi/512
   cos[287]  =  13'b1111001111101;     //287pi/512
   sin[288]  =  13'b1100000100111;     //288pi/512
   cos[288]  =  13'b1111001110000;     //288pi/512
   sin[289]  =  13'b1100000101010;     //289pi/512
   cos[289]  =  13'b1111001100100;     //289pi/512
   sin[290]  =  13'b1100000101100;     //290pi/512
   cos[290]  =  13'b1111001011000;     //290pi/512
   sin[291]  =  13'b1100000101111;     //291pi/512
   cos[291]  =  13'b1111001001100;     //291pi/512
   sin[292]  =  13'b1100000110010;     //292pi/512
   cos[292]  =  13'b1111000111111;     //292pi/512
   sin[293]  =  13'b1100000110101;     //293pi/512
   cos[293]  =  13'b1111000110011;     //293pi/512
   sin[294]  =  13'b1100000110111;     //294pi/512
   cos[294]  =  13'b1111000100111;     //294pi/512
   sin[295]  =  13'b1100000111010;     //295pi/512
   cos[295]  =  13'b1111000011011;     //295pi/512
   sin[296]  =  13'b1100000111101;     //296pi/512
   cos[296]  =  13'b1111000001110;     //296pi/512
   sin[297]  =  13'b1100001000000;     //297pi/512
   cos[297]  =  13'b1111000000010;     //297pi/512
   sin[298]  =  13'b1100001000100;     //298pi/512
   cos[298]  =  13'b1110111110110;     //298pi/512
   sin[299]  =  13'b1100001000111;     //299pi/512
   cos[299]  =  13'b1110111101010;     //299pi/512
   sin[300]  =  13'b1100001001010;     //300pi/512
   cos[300]  =  13'b1110111011110;     //300pi/512
   sin[301]  =  13'b1100001001110;     //301pi/512
   cos[301]  =  13'b1110111010010;     //301pi/512
   sin[302]  =  13'b1100001010001;     //302pi/512
   cos[302]  =  13'b1110111000110;     //302pi/512
   sin[303]  =  13'b1100001010101;     //303pi/512
   cos[303]  =  13'b1110110111010;     //303pi/512
   sin[304]  =  13'b1100001011000;     //304pi/512
   cos[304]  =  13'b1110110101101;     //304pi/512
   sin[305]  =  13'b1100001011100;     //305pi/512
   cos[305]  =  13'b1110110100001;     //305pi/512
   sin[306]  =  13'b1100001100000;     //306pi/512
   cos[306]  =  13'b1110110010101;     //306pi/512
   sin[307]  =  13'b1100001100011;     //307pi/512
   cos[307]  =  13'b1110110001010;     //307pi/512
   sin[308]  =  13'b1100001100111;     //308pi/512
   cos[308]  =  13'b1110101111110;     //308pi/512
   sin[309]  =  13'b1100001101011;     //309pi/512
   cos[309]  =  13'b1110101110010;     //309pi/512
   sin[310]  =  13'b1100001101111;     //310pi/512
   cos[310]  =  13'b1110101100110;     //310pi/512
   sin[311]  =  13'b1100001110100;     //311pi/512
   cos[311]  =  13'b1110101011010;     //311pi/512
   sin[312]  =  13'b1100001111000;     //312pi/512
   cos[312]  =  13'b1110101001110;     //312pi/512
   sin[313]  =  13'b1100001111100;     //313pi/512
   cos[313]  =  13'b1110101000010;     //313pi/512
   sin[314]  =  13'b1100010000000;     //314pi/512
   cos[314]  =  13'b1110100110110;     //314pi/512
   sin[315]  =  13'b1100010000101;     //315pi/512
   cos[315]  =  13'b1110100101011;     //315pi/512
   sin[316]  =  13'b1100010001001;     //316pi/512
   cos[316]  =  13'b1110100011111;     //316pi/512
   sin[317]  =  13'b1100010001110;     //317pi/512
   cos[317]  =  13'b1110100010011;     //317pi/512
   sin[318]  =  13'b1100010010010;     //318pi/512
   cos[318]  =  13'b1110100001000;     //318pi/512
   sin[319]  =  13'b1100010010111;     //319pi/512
   cos[319]  =  13'b1110011111100;     //319pi/512
   sin[320]  =  13'b1100010011100;     //320pi/512
   cos[320]  =  13'b1110011110000;     //320pi/512
   sin[321]  =  13'b1100010100001;     //321pi/512
   cos[321]  =  13'b1110011100101;     //321pi/512
   sin[322]  =  13'b1100010100110;     //322pi/512
   cos[322]  =  13'b1110011011001;     //322pi/512
   sin[323]  =  13'b1100010101011;     //323pi/512
   cos[323]  =  13'b1110011001110;     //323pi/512
   sin[324]  =  13'b1100010110000;     //324pi/512
   cos[324]  =  13'b1110011000010;     //324pi/512
   sin[325]  =  13'b1100010110101;     //325pi/512
   cos[325]  =  13'b1110010110111;     //325pi/512
   sin[326]  =  13'b1100010111010;     //326pi/512
   cos[326]  =  13'b1110010101011;     //326pi/512
   sin[327]  =  13'b1100010111111;     //327pi/512
   cos[327]  =  13'b1110010100000;     //327pi/512
   sin[328]  =  13'b1100011000101;     //328pi/512
   cos[328]  =  13'b1110010010100;     //328pi/512
   sin[329]  =  13'b1100011001010;     //329pi/512
   cos[329]  =  13'b1110010001001;     //329pi/512
   sin[330]  =  13'b1100011010000;     //330pi/512
   cos[330]  =  13'b1110001111110;     //330pi/512
   sin[331]  =  13'b1100011010101;     //331pi/512
   cos[331]  =  13'b1110001110010;     //331pi/512
   sin[332]  =  13'b1100011011011;     //332pi/512
   cos[332]  =  13'b1110001100111;     //332pi/512
   sin[333]  =  13'b1100011100000;     //333pi/512
   cos[333]  =  13'b1110001011100;     //333pi/512
   sin[334]  =  13'b1100011100110;     //334pi/512
   cos[334]  =  13'b1110001010001;     //334pi/512
   sin[335]  =  13'b1100011101100;     //335pi/512
   cos[335]  =  13'b1110001000110;     //335pi/512
   sin[336]  =  13'b1100011110010;     //336pi/512
   cos[336]  =  13'b1110000111011;     //336pi/512
   sin[337]  =  13'b1100011111000;     //337pi/512
   cos[337]  =  13'b1110000110000;     //337pi/512
   sin[338]  =  13'b1100011111110;     //338pi/512
   cos[338]  =  13'b1110000100100;     //338pi/512
   sin[339]  =  13'b1100100000100;     //339pi/512
   cos[339]  =  13'b1110000011001;     //339pi/512
   sin[340]  =  13'b1100100001010;     //340pi/512
   cos[340]  =  13'b1110000001111;     //340pi/512
   sin[341]  =  13'b1100100010000;     //341pi/512
   cos[341]  =  13'b1110000000100;     //341pi/512
   sin[342]  =  13'b1100100010111;     //342pi/512
   cos[342]  =  13'b1101111111001;     //342pi/512
   sin[343]  =  13'b1100100011101;     //343pi/512
   cos[343]  =  13'b1101111101110;     //343pi/512
   sin[344]  =  13'b1100100100011;     //344pi/512
   cos[344]  =  13'b1101111100011;     //344pi/512
   sin[345]  =  13'b1100100101010;     //345pi/512
   cos[345]  =  13'b1101111011000;     //345pi/512
   sin[346]  =  13'b1100100110000;     //346pi/512
   cos[346]  =  13'b1101111001110;     //346pi/512
   sin[347]  =  13'b1100100110111;     //347pi/512
   cos[347]  =  13'b1101111000011;     //347pi/512
   sin[348]  =  13'b1100100111110;     //348pi/512
   cos[348]  =  13'b1101110111000;     //348pi/512
   sin[349]  =  13'b1100101000100;     //349pi/512
   cos[349]  =  13'b1101110101110;     //349pi/512
   sin[350]  =  13'b1100101001011;     //350pi/512
   cos[350]  =  13'b1101110100011;     //350pi/512
   sin[351]  =  13'b1100101010010;     //351pi/512
   cos[351]  =  13'b1101110011001;     //351pi/512
   sin[352]  =  13'b1100101011001;     //352pi/512
   cos[352]  =  13'b1101110001110;     //352pi/512
   sin[353]  =  13'b1100101100000;     //353pi/512
   cos[353]  =  13'b1101110000100;     //353pi/512
   sin[354]  =  13'b1100101100111;     //354pi/512
   cos[354]  =  13'b1101101111001;     //354pi/512
   sin[355]  =  13'b1100101101110;     //355pi/512
   cos[355]  =  13'b1101101101111;     //355pi/512
   sin[356]  =  13'b1100101110110;     //356pi/512
   cos[356]  =  13'b1101101100101;     //356pi/512
   sin[357]  =  13'b1100101111101;     //357pi/512
   cos[357]  =  13'b1101101011010;     //357pi/512
   sin[358]  =  13'b1100110000100;     //358pi/512
   cos[358]  =  13'b1101101010000;     //358pi/512
   sin[359]  =  13'b1100110001100;     //359pi/512
   cos[359]  =  13'b1101101000110;     //359pi/512
   sin[360]  =  13'b1100110010011;     //360pi/512
   cos[360]  =  13'b1101100111100;     //360pi/512
   sin[361]  =  13'b1100110011011;     //361pi/512
   cos[361]  =  13'b1101100110010;     //361pi/512
   sin[362]  =  13'b1100110100010;     //362pi/512
   cos[362]  =  13'b1101100101000;     //362pi/512
   sin[363]  =  13'b1100110101010;     //363pi/512
   cos[363]  =  13'b1101100011110;     //363pi/512
   sin[364]  =  13'b1100110110001;     //364pi/512
   cos[364]  =  13'b1101100010100;     //364pi/512
   sin[365]  =  13'b1100110111001;     //365pi/512
   cos[365]  =  13'b1101100001010;     //365pi/512
   sin[366]  =  13'b1100111000001;     //366pi/512
   cos[366]  =  13'b1101100000000;     //366pi/512
   sin[367]  =  13'b1100111001001;     //367pi/512
   cos[367]  =  13'b1101011110111;     //367pi/512
   sin[368]  =  13'b1100111010001;     //368pi/512
   cos[368]  =  13'b1101011101101;     //368pi/512
   sin[369]  =  13'b1100111011001;     //369pi/512
   cos[369]  =  13'b1101011100011;     //369pi/512
   sin[370]  =  13'b1100111100001;     //370pi/512
   cos[370]  =  13'b1101011011001;     //370pi/512
   sin[371]  =  13'b1100111101001;     //371pi/512
   cos[371]  =  13'b1101011010000;     //371pi/512
   sin[372]  =  13'b1100111110001;     //372pi/512
   cos[372]  =  13'b1101011000110;     //372pi/512
   sin[373]  =  13'b1100111111001;     //373pi/512
   cos[373]  =  13'b1101010111101;     //373pi/512
   sin[374]  =  13'b1101000000010;     //374pi/512
   cos[374]  =  13'b1101010110011;     //374pi/512
   sin[375]  =  13'b1101000001010;     //375pi/512
   cos[375]  =  13'b1101010101010;     //375pi/512
   sin[376]  =  13'b1101000010011;     //376pi/512
   cos[376]  =  13'b1101010100001;     //376pi/512
   sin[377]  =  13'b1101000011011;     //377pi/512
   cos[377]  =  13'b1101010010111;     //377pi/512
   sin[378]  =  13'b1101000100100;     //378pi/512
   cos[378]  =  13'b1101010001110;     //378pi/512
   sin[379]  =  13'b1101000101100;     //379pi/512
   cos[379]  =  13'b1101010000101;     //379pi/512
   sin[380]  =  13'b1101000110101;     //380pi/512
   cos[380]  =  13'b1101001111100;     //380pi/512
   sin[381]  =  13'b1101000111101;     //381pi/512
   cos[381]  =  13'b1101001110011;     //381pi/512
   sin[382]  =  13'b1101001000110;     //382pi/512
   cos[382]  =  13'b1101001101010;     //382pi/512
   sin[383]  =  13'b1101001001111;     //383pi/512
   cos[383]  =  13'b1101001100001;     //383pi/512
   sin[384]  =  13'b1101001011000;     //384pi/512
   cos[384]  =  13'b1101001011000;     //384pi/512
   sin[385]  =  13'b1101001100001;     //385pi/512
   cos[385]  =  13'b1101001001111;     //385pi/512
   sin[386]  =  13'b1101001101010;     //386pi/512
   cos[386]  =  13'b1101001000110;     //386pi/512
   sin[387]  =  13'b1101001110011;     //387pi/512
   cos[387]  =  13'b1101000111101;     //387pi/512
   sin[388]  =  13'b1101001111100;     //388pi/512
   cos[388]  =  13'b1101000110101;     //388pi/512
   sin[389]  =  13'b1101010000101;     //389pi/512
   cos[389]  =  13'b1101000101100;     //389pi/512
   sin[390]  =  13'b1101010001110;     //390pi/512
   cos[390]  =  13'b1101000100100;     //390pi/512
   sin[391]  =  13'b1101010010111;     //391pi/512
   cos[391]  =  13'b1101000011011;     //391pi/512
   sin[392]  =  13'b1101010100001;     //392pi/512
   cos[392]  =  13'b1101000010011;     //392pi/512
   sin[393]  =  13'b1101010101010;     //393pi/512
   cos[393]  =  13'b1101000001010;     //393pi/512
   sin[394]  =  13'b1101010110011;     //394pi/512
   cos[394]  =  13'b1101000000010;     //394pi/512
   sin[395]  =  13'b1101010111101;     //395pi/512
   cos[395]  =  13'b1100111111001;     //395pi/512
   sin[396]  =  13'b1101011000110;     //396pi/512
   cos[396]  =  13'b1100111110001;     //396pi/512
   sin[397]  =  13'b1101011010000;     //397pi/512
   cos[397]  =  13'b1100111101001;     //397pi/512
   sin[398]  =  13'b1101011011001;     //398pi/512
   cos[398]  =  13'b1100111100001;     //398pi/512
   sin[399]  =  13'b1101011100011;     //399pi/512
   cos[399]  =  13'b1100111011001;     //399pi/512
   sin[400]  =  13'b1101011101101;     //400pi/512
   cos[400]  =  13'b1100111010001;     //400pi/512
   sin[401]  =  13'b1101011110111;     //401pi/512
   cos[401]  =  13'b1100111001001;     //401pi/512
   sin[402]  =  13'b1101100000000;     //402pi/512
   cos[402]  =  13'b1100111000001;     //402pi/512
   sin[403]  =  13'b1101100001010;     //403pi/512
   cos[403]  =  13'b1100110111001;     //403pi/512
   sin[404]  =  13'b1101100010100;     //404pi/512
   cos[404]  =  13'b1100110110001;     //404pi/512
   sin[405]  =  13'b1101100011110;     //405pi/512
   cos[405]  =  13'b1100110101010;     //405pi/512
   sin[406]  =  13'b1101100101000;     //406pi/512
   cos[406]  =  13'b1100110100010;     //406pi/512
   sin[407]  =  13'b1101100110010;     //407pi/512
   cos[407]  =  13'b1100110011011;     //407pi/512
   sin[408]  =  13'b1101100111100;     //408pi/512
   cos[408]  =  13'b1100110010011;     //408pi/512
   sin[409]  =  13'b1101101000110;     //409pi/512
   cos[409]  =  13'b1100110001100;     //409pi/512
   sin[410]  =  13'b1101101010000;     //410pi/512
   cos[410]  =  13'b1100110000100;     //410pi/512
   sin[411]  =  13'b1101101011010;     //411pi/512
   cos[411]  =  13'b1100101111101;     //411pi/512
   sin[412]  =  13'b1101101100101;     //412pi/512
   cos[412]  =  13'b1100101110110;     //412pi/512
   sin[413]  =  13'b1101101101111;     //413pi/512
   cos[413]  =  13'b1100101101110;     //413pi/512
   sin[414]  =  13'b1101101111001;     //414pi/512
   cos[414]  =  13'b1100101100111;     //414pi/512
   sin[415]  =  13'b1101110000100;     //415pi/512
   cos[415]  =  13'b1100101100000;     //415pi/512
   sin[416]  =  13'b1101110001110;     //416pi/512
   cos[416]  =  13'b1100101011001;     //416pi/512
   sin[417]  =  13'b1101110011001;     //417pi/512
   cos[417]  =  13'b1100101010010;     //417pi/512
   sin[418]  =  13'b1101110100011;     //418pi/512
   cos[418]  =  13'b1100101001011;     //418pi/512
   sin[419]  =  13'b1101110101110;     //419pi/512
   cos[419]  =  13'b1100101000100;     //419pi/512
   sin[420]  =  13'b1101110111000;     //420pi/512
   cos[420]  =  13'b1100100111110;     //420pi/512
   sin[421]  =  13'b1101111000011;     //421pi/512
   cos[421]  =  13'b1100100110111;     //421pi/512
   sin[422]  =  13'b1101111001110;     //422pi/512
   cos[422]  =  13'b1100100110000;     //422pi/512
   sin[423]  =  13'b1101111011000;     //423pi/512
   cos[423]  =  13'b1100100101010;     //423pi/512
   sin[424]  =  13'b1101111100011;     //424pi/512
   cos[424]  =  13'b1100100100011;     //424pi/512
   sin[425]  =  13'b1101111101110;     //425pi/512
   cos[425]  =  13'b1100100011101;     //425pi/512
   sin[426]  =  13'b1101111111001;     //426pi/512
   cos[426]  =  13'b1100100010111;     //426pi/512
   sin[427]  =  13'b1110000000100;     //427pi/512
   cos[427]  =  13'b1100100010000;     //427pi/512
   sin[428]  =  13'b1110000001111;     //428pi/512
   cos[428]  =  13'b1100100001010;     //428pi/512
   sin[429]  =  13'b1110000011001;     //429pi/512
   cos[429]  =  13'b1100100000100;     //429pi/512
   sin[430]  =  13'b1110000100100;     //430pi/512
   cos[430]  =  13'b1100011111110;     //430pi/512
   sin[431]  =  13'b1110000110000;     //431pi/512
   cos[431]  =  13'b1100011111000;     //431pi/512
   sin[432]  =  13'b1110000111011;     //432pi/512
   cos[432]  =  13'b1100011110010;     //432pi/512
   sin[433]  =  13'b1110001000110;     //433pi/512
   cos[433]  =  13'b1100011101100;     //433pi/512
   sin[434]  =  13'b1110001010001;     //434pi/512
   cos[434]  =  13'b1100011100110;     //434pi/512
   sin[435]  =  13'b1110001011100;     //435pi/512
   cos[435]  =  13'b1100011100000;     //435pi/512
   sin[436]  =  13'b1110001100111;     //436pi/512
   cos[436]  =  13'b1100011011011;     //436pi/512
   sin[437]  =  13'b1110001110010;     //437pi/512
   cos[437]  =  13'b1100011010101;     //437pi/512
   sin[438]  =  13'b1110001111110;     //438pi/512
   cos[438]  =  13'b1100011010000;     //438pi/512
   sin[439]  =  13'b1110010001001;     //439pi/512
   cos[439]  =  13'b1100011001010;     //439pi/512
   sin[440]  =  13'b1110010010100;     //440pi/512
   cos[440]  =  13'b1100011000101;     //440pi/512
   sin[441]  =  13'b1110010100000;     //441pi/512
   cos[441]  =  13'b1100010111111;     //441pi/512
   sin[442]  =  13'b1110010101011;     //442pi/512
   cos[442]  =  13'b1100010111010;     //442pi/512
   sin[443]  =  13'b1110010110111;     //443pi/512
   cos[443]  =  13'b1100010110101;     //443pi/512
   sin[444]  =  13'b1110011000010;     //444pi/512
   cos[444]  =  13'b1100010110000;     //444pi/512
   sin[445]  =  13'b1110011001110;     //445pi/512
   cos[445]  =  13'b1100010101011;     //445pi/512
   sin[446]  =  13'b1110011011001;     //446pi/512
   cos[446]  =  13'b1100010100110;     //446pi/512
   sin[447]  =  13'b1110011100101;     //447pi/512
   cos[447]  =  13'b1100010100001;     //447pi/512
   sin[448]  =  13'b1110011110000;     //448pi/512
   cos[448]  =  13'b1100010011100;     //448pi/512
   sin[449]  =  13'b1110011111100;     //449pi/512
   cos[449]  =  13'b1100010010111;     //449pi/512
   sin[450]  =  13'b1110100001000;     //450pi/512
   cos[450]  =  13'b1100010010010;     //450pi/512
   sin[451]  =  13'b1110100010011;     //451pi/512
   cos[451]  =  13'b1100010001110;     //451pi/512
   sin[452]  =  13'b1110100011111;     //452pi/512
   cos[452]  =  13'b1100010001001;     //452pi/512
   sin[453]  =  13'b1110100101011;     //453pi/512
   cos[453]  =  13'b1100010000101;     //453pi/512
   sin[454]  =  13'b1110100110110;     //454pi/512
   cos[454]  =  13'b1100010000000;     //454pi/512
   sin[455]  =  13'b1110101000010;     //455pi/512
   cos[455]  =  13'b1100001111100;     //455pi/512
   sin[456]  =  13'b1110101001110;     //456pi/512
   cos[456]  =  13'b1100001111000;     //456pi/512
   sin[457]  =  13'b1110101011010;     //457pi/512
   cos[457]  =  13'b1100001110100;     //457pi/512
   sin[458]  =  13'b1110101100110;     //458pi/512
   cos[458]  =  13'b1100001101111;     //458pi/512
   sin[459]  =  13'b1110101110010;     //459pi/512
   cos[459]  =  13'b1100001101011;     //459pi/512
   sin[460]  =  13'b1110101111110;     //460pi/512
   cos[460]  =  13'b1100001100111;     //460pi/512
   sin[461]  =  13'b1110110001010;     //461pi/512
   cos[461]  =  13'b1100001100011;     //461pi/512
   sin[462]  =  13'b1110110010101;     //462pi/512
   cos[462]  =  13'b1100001100000;     //462pi/512
   sin[463]  =  13'b1110110100001;     //463pi/512
   cos[463]  =  13'b1100001011100;     //463pi/512
   sin[464]  =  13'b1110110101101;     //464pi/512
   cos[464]  =  13'b1100001011000;     //464pi/512
   sin[465]  =  13'b1110110111010;     //465pi/512
   cos[465]  =  13'b1100001010101;     //465pi/512
   sin[466]  =  13'b1110111000110;     //466pi/512
   cos[466]  =  13'b1100001010001;     //466pi/512
   sin[467]  =  13'b1110111010010;     //467pi/512
   cos[467]  =  13'b1100001001110;     //467pi/512
   sin[468]  =  13'b1110111011110;     //468pi/512
   cos[468]  =  13'b1100001001010;     //468pi/512
   sin[469]  =  13'b1110111101010;     //469pi/512
   cos[469]  =  13'b1100001000111;     //469pi/512
   sin[470]  =  13'b1110111110110;     //470pi/512
   cos[470]  =  13'b1100001000100;     //470pi/512
   sin[471]  =  13'b1111000000010;     //471pi/512
   cos[471]  =  13'b1100001000000;     //471pi/512
   sin[472]  =  13'b1111000001110;     //472pi/512
   cos[472]  =  13'b1100000111101;     //472pi/512
   sin[473]  =  13'b1111000011011;     //473pi/512
   cos[473]  =  13'b1100000111010;     //473pi/512
   sin[474]  =  13'b1111000100111;     //474pi/512
   cos[474]  =  13'b1100000110111;     //474pi/512
   sin[475]  =  13'b1111000110011;     //475pi/512
   cos[475]  =  13'b1100000110101;     //475pi/512
   sin[476]  =  13'b1111000111111;     //476pi/512
   cos[476]  =  13'b1100000110010;     //476pi/512
   sin[477]  =  13'b1111001001100;     //477pi/512
   cos[477]  =  13'b1100000101111;     //477pi/512
   sin[478]  =  13'b1111001011000;     //478pi/512
   cos[478]  =  13'b1100000101100;     //478pi/512
   sin[479]  =  13'b1111001100100;     //479pi/512
   cos[479]  =  13'b1100000101010;     //479pi/512
   sin[480]  =  13'b1111001110000;     //480pi/512
   cos[480]  =  13'b1100000100111;     //480pi/512
   sin[481]  =  13'b1111001111101;     //481pi/512
   cos[481]  =  13'b1100000100101;     //481pi/512
   sin[482]  =  13'b1111010001001;     //482pi/512
   cos[482]  =  13'b1100000100011;     //482pi/512
   sin[483]  =  13'b1111010010101;     //483pi/512
   cos[483]  =  13'b1100000100000;     //483pi/512
   sin[484]  =  13'b1111010100010;     //484pi/512
   cos[484]  =  13'b1100000011110;     //484pi/512
   sin[485]  =  13'b1111010101110;     //485pi/512
   cos[485]  =  13'b1100000011100;     //485pi/512
   sin[486]  =  13'b1111010111011;     //486pi/512
   cos[486]  =  13'b1100000011010;     //486pi/512
   sin[487]  =  13'b1111011000111;     //487pi/512
   cos[487]  =  13'b1100000011000;     //487pi/512
   sin[488]  =  13'b1111011010011;     //488pi/512
   cos[488]  =  13'b1100000010110;     //488pi/512
   sin[489]  =  13'b1111011100000;     //489pi/512
   cos[489]  =  13'b1100000010100;     //489pi/512
   sin[490]  =  13'b1111011101100;     //490pi/512
   cos[490]  =  13'b1100000010011;     //490pi/512
   sin[491]  =  13'b1111011111001;     //491pi/512
   cos[491]  =  13'b1100000010001;     //491pi/512
   sin[492]  =  13'b1111100000101;     //492pi/512
   cos[492]  =  13'b1100000001111;     //492pi/512
   sin[493]  =  13'b1111100010010;     //493pi/512
   cos[493]  =  13'b1100000001110;     //493pi/512
   sin[494]  =  13'b1111100011110;     //494pi/512
   cos[494]  =  13'b1100000001100;     //494pi/512
   sin[495]  =  13'b1111100101011;     //495pi/512
   cos[495]  =  13'b1100000001011;     //495pi/512
   sin[496]  =  13'b1111100110111;     //496pi/512
   cos[496]  =  13'b1100000001010;     //496pi/512
   sin[497]  =  13'b1111101000100;     //497pi/512
   cos[497]  =  13'b1100000001001;     //497pi/512
   sin[498]  =  13'b1111101010000;     //498pi/512
   cos[498]  =  13'b1100000001000;     //498pi/512
   sin[499]  =  13'b1111101011101;     //499pi/512
   cos[499]  =  13'b1100000000111;     //499pi/512
   sin[500]  =  13'b1111101101001;     //500pi/512
   cos[500]  =  13'b1100000000110;     //500pi/512
   sin[501]  =  13'b1111101110110;     //501pi/512
   cos[501]  =  13'b1100000000101;     //501pi/512
   sin[502]  =  13'b1111110000010;     //502pi/512
   cos[502]  =  13'b1100000000100;     //502pi/512
   sin[503]  =  13'b1111110001111;     //503pi/512
   cos[503]  =  13'b1100000000011;     //503pi/512
   sin[504]  =  13'b1111110011100;     //504pi/512
   cos[504]  =  13'b1100000000010;     //504pi/512
   sin[505]  =  13'b1111110101000;     //505pi/512
   cos[505]  =  13'b1100000000010;     //505pi/512
   sin[506]  =  13'b1111110110101;     //506pi/512
   cos[506]  =  13'b1100000000001;     //506pi/512
   sin[507]  =  13'b1111111000001;     //507pi/512
   cos[507]  =  13'b1100000000001;     //507pi/512
   sin[508]  =  13'b1111111001110;     //508pi/512
   cos[508]  =  13'b1100000000001;     //508pi/512
   sin[509]  =  13'b1111111011010;     //509pi/512
   cos[509]  =  13'b1100000000000;     //509pi/512
   sin[510]  =  13'b1111111100111;     //510pi/512
   cos[510]  =  13'b1100000000000;     //510pi/512
   sin[511]  =  13'b1111111110011;     //511pi/512
   cos[511]  =  13'b1100000000000;     //511pi/512
end
endmodule
