module  TWIDLE_9_bit  #(parameter SIZE = 10, word_length_tw = 9) (
    input            clk,
    input            en_rd,
    input   [10:0]   rd_ptr_angle,
    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );
reg signed [word_length_tw-1:0]  cos  [511:0];
reg signed [word_length_tw-1:0]  sin  [511:0];
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd) begin
                  cos_data           <= cos   [rd_ptr_angle];
                  sin_data           <= sin   [rd_ptr_angle];
             end 
        end
initial begin
   sin[0]  =  9'b000000000;     //0pi/512
   cos[0]  =  9'b010000000;     //0pi/512
   sin[1]  =  9'b111111111;     //1pi/512
   cos[1]  =  9'b001111111;     //1pi/512
   sin[2]  =  9'b111111110;     //2pi/512
   cos[2]  =  9'b001111111;     //2pi/512
   sin[3]  =  9'b111111110;     //3pi/512
   cos[3]  =  9'b001111111;     //3pi/512
   sin[4]  =  9'b111111101;     //4pi/512
   cos[4]  =  9'b001111111;     //4pi/512
   sin[5]  =  9'b111111100;     //5pi/512
   cos[5]  =  9'b001111111;     //5pi/512
   sin[6]  =  9'b111111011;     //6pi/512
   cos[6]  =  9'b001111111;     //6pi/512
   sin[7]  =  9'b111111011;     //7pi/512
   cos[7]  =  9'b001111111;     //7pi/512
   sin[8]  =  9'b111111010;     //8pi/512
   cos[8]  =  9'b001111111;     //8pi/512
   sin[9]  =  9'b111111001;     //9pi/512
   cos[9]  =  9'b001111111;     //9pi/512
   sin[10]  =  9'b111111000;     //10pi/512
   cos[10]  =  9'b001111111;     //10pi/512
   sin[11]  =  9'b111110111;     //11pi/512
   cos[11]  =  9'b001111111;     //11pi/512
   sin[12]  =  9'b111110111;     //12pi/512
   cos[12]  =  9'b001111111;     //12pi/512
   sin[13]  =  9'b111110110;     //13pi/512
   cos[13]  =  9'b001111111;     //13pi/512
   sin[14]  =  9'b111110101;     //14pi/512
   cos[14]  =  9'b001111111;     //14pi/512
   sin[15]  =  9'b111110100;     //15pi/512
   cos[15]  =  9'b001111111;     //15pi/512
   sin[16]  =  9'b111110011;     //16pi/512
   cos[16]  =  9'b001111111;     //16pi/512
   sin[17]  =  9'b111110011;     //17pi/512
   cos[17]  =  9'b001111111;     //17pi/512
   sin[18]  =  9'b111110010;     //18pi/512
   cos[18]  =  9'b001111111;     //18pi/512
   sin[19]  =  9'b111110001;     //19pi/512
   cos[19]  =  9'b001111111;     //19pi/512
   sin[20]  =  9'b111110000;     //20pi/512
   cos[20]  =  9'b001111111;     //20pi/512
   sin[21]  =  9'b111110000;     //21pi/512
   cos[21]  =  9'b001111110;     //21pi/512
   sin[22]  =  9'b111101111;     //22pi/512
   cos[22]  =  9'b001111110;     //22pi/512
   sin[23]  =  9'b111101110;     //23pi/512
   cos[23]  =  9'b001111110;     //23pi/512
   sin[24]  =  9'b111101101;     //24pi/512
   cos[24]  =  9'b001111110;     //24pi/512
   sin[25]  =  9'b111101100;     //25pi/512
   cos[25]  =  9'b001111110;     //25pi/512
   sin[26]  =  9'b111101100;     //26pi/512
   cos[26]  =  9'b001111110;     //26pi/512
   sin[27]  =  9'b111101011;     //27pi/512
   cos[27]  =  9'b001111110;     //27pi/512
   sin[28]  =  9'b111101010;     //28pi/512
   cos[28]  =  9'b001111110;     //28pi/512
   sin[29]  =  9'b111101001;     //29pi/512
   cos[29]  =  9'b001111101;     //29pi/512
   sin[30]  =  9'b111101001;     //30pi/512
   cos[30]  =  9'b001111101;     //30pi/512
   sin[31]  =  9'b111101000;     //31pi/512
   cos[31]  =  9'b001111101;     //31pi/512
   sin[32]  =  9'b111100111;     //32pi/512
   cos[32]  =  9'b001111101;     //32pi/512
   sin[33]  =  9'b111100110;     //33pi/512
   cos[33]  =  9'b001111101;     //33pi/512
   sin[34]  =  9'b111100101;     //34pi/512
   cos[34]  =  9'b001111101;     //34pi/512
   sin[35]  =  9'b111100101;     //35pi/512
   cos[35]  =  9'b001111101;     //35pi/512
   sin[36]  =  9'b111100100;     //36pi/512
   cos[36]  =  9'b001111100;     //36pi/512
   sin[37]  =  9'b111100011;     //37pi/512
   cos[37]  =  9'b001111100;     //37pi/512
   sin[38]  =  9'b111100010;     //38pi/512
   cos[38]  =  9'b001111100;     //38pi/512
   sin[39]  =  9'b111100010;     //39pi/512
   cos[39]  =  9'b001111100;     //39pi/512
   sin[40]  =  9'b111100001;     //40pi/512
   cos[40]  =  9'b001111100;     //40pi/512
   sin[41]  =  9'b111100000;     //41pi/512
   cos[41]  =  9'b001111011;     //41pi/512
   sin[42]  =  9'b111011111;     //42pi/512
   cos[42]  =  9'b001111011;     //42pi/512
   sin[43]  =  9'b111011111;     //43pi/512
   cos[43]  =  9'b001111011;     //43pi/512
   sin[44]  =  9'b111011110;     //44pi/512
   cos[44]  =  9'b001111011;     //44pi/512
   sin[45]  =  9'b111011101;     //45pi/512
   cos[45]  =  9'b001111011;     //45pi/512
   sin[46]  =  9'b111011100;     //46pi/512
   cos[46]  =  9'b001111010;     //46pi/512
   sin[47]  =  9'b111011100;     //47pi/512
   cos[47]  =  9'b001111010;     //47pi/512
   sin[48]  =  9'b111011011;     //48pi/512
   cos[48]  =  9'b001111010;     //48pi/512
   sin[49]  =  9'b111011010;     //49pi/512
   cos[49]  =  9'b001111010;     //49pi/512
   sin[50]  =  9'b111011001;     //50pi/512
   cos[50]  =  9'b001111010;     //50pi/512
   sin[51]  =  9'b111011001;     //51pi/512
   cos[51]  =  9'b001111001;     //51pi/512
   sin[52]  =  9'b111011000;     //52pi/512
   cos[52]  =  9'b001111001;     //52pi/512
   sin[53]  =  9'b111010111;     //53pi/512
   cos[53]  =  9'b001111001;     //53pi/512
   sin[54]  =  9'b111010110;     //54pi/512
   cos[54]  =  9'b001111001;     //54pi/512
   sin[55]  =  9'b111010110;     //55pi/512
   cos[55]  =  9'b001111000;     //55pi/512
   sin[56]  =  9'b111010101;     //56pi/512
   cos[56]  =  9'b001111000;     //56pi/512
   sin[57]  =  9'b111010100;     //57pi/512
   cos[57]  =  9'b001111000;     //57pi/512
   sin[58]  =  9'b111010011;     //58pi/512
   cos[58]  =  9'b001110111;     //58pi/512
   sin[59]  =  9'b111010011;     //59pi/512
   cos[59]  =  9'b001110111;     //59pi/512
   sin[60]  =  9'b111010010;     //60pi/512
   cos[60]  =  9'b001110111;     //60pi/512
   sin[61]  =  9'b111010001;     //61pi/512
   cos[61]  =  9'b001110111;     //61pi/512
   sin[62]  =  9'b111010000;     //62pi/512
   cos[62]  =  9'b001110110;     //62pi/512
   sin[63]  =  9'b111010000;     //63pi/512
   cos[63]  =  9'b001110110;     //63pi/512
   sin[64]  =  9'b111001111;     //64pi/512
   cos[64]  =  9'b001110110;     //64pi/512
   sin[65]  =  9'b111001110;     //65pi/512
   cos[65]  =  9'b001110101;     //65pi/512
   sin[66]  =  9'b111001110;     //66pi/512
   cos[66]  =  9'b001110101;     //66pi/512
   sin[67]  =  9'b111001101;     //67pi/512
   cos[67]  =  9'b001110101;     //67pi/512
   sin[68]  =  9'b111001100;     //68pi/512
   cos[68]  =  9'b001110101;     //68pi/512
   sin[69]  =  9'b111001011;     //69pi/512
   cos[69]  =  9'b001110100;     //69pi/512
   sin[70]  =  9'b111001011;     //70pi/512
   cos[70]  =  9'b001110100;     //70pi/512
   sin[71]  =  9'b111001010;     //71pi/512
   cos[71]  =  9'b001110100;     //71pi/512
   sin[72]  =  9'b111001001;     //72pi/512
   cos[72]  =  9'b001110011;     //72pi/512
   sin[73]  =  9'b111001001;     //73pi/512
   cos[73]  =  9'b001110011;     //73pi/512
   sin[74]  =  9'b111001000;     //74pi/512
   cos[74]  =  9'b001110011;     //74pi/512
   sin[75]  =  9'b111000111;     //75pi/512
   cos[75]  =  9'b001110010;     //75pi/512
   sin[76]  =  9'b111000110;     //76pi/512
   cos[76]  =  9'b001110010;     //76pi/512
   sin[77]  =  9'b111000110;     //77pi/512
   cos[77]  =  9'b001110001;     //77pi/512
   sin[78]  =  9'b111000101;     //78pi/512
   cos[78]  =  9'b001110001;     //78pi/512
   sin[79]  =  9'b111000100;     //79pi/512
   cos[79]  =  9'b001110001;     //79pi/512
   sin[80]  =  9'b111000100;     //80pi/512
   cos[80]  =  9'b001110000;     //80pi/512
   sin[81]  =  9'b111000011;     //81pi/512
   cos[81]  =  9'b001110000;     //81pi/512
   sin[82]  =  9'b111000010;     //82pi/512
   cos[82]  =  9'b001110000;     //82pi/512
   sin[83]  =  9'b111000010;     //83pi/512
   cos[83]  =  9'b001101111;     //83pi/512
   sin[84]  =  9'b111000001;     //84pi/512
   cos[84]  =  9'b001101111;     //84pi/512
   sin[85]  =  9'b111000000;     //85pi/512
   cos[85]  =  9'b001101110;     //85pi/512
   sin[86]  =  9'b111000000;     //86pi/512
   cos[86]  =  9'b001101110;     //86pi/512
   sin[87]  =  9'b110111111;     //87pi/512
   cos[87]  =  9'b001101110;     //87pi/512
   sin[88]  =  9'b110111110;     //88pi/512
   cos[88]  =  9'b001101101;     //88pi/512
   sin[89]  =  9'b110111110;     //89pi/512
   cos[89]  =  9'b001101101;     //89pi/512
   sin[90]  =  9'b110111101;     //90pi/512
   cos[90]  =  9'b001101100;     //90pi/512
   sin[91]  =  9'b110111100;     //91pi/512
   cos[91]  =  9'b001101100;     //91pi/512
   sin[92]  =  9'b110111100;     //92pi/512
   cos[92]  =  9'b001101100;     //92pi/512
   sin[93]  =  9'b110111011;     //93pi/512
   cos[93]  =  9'b001101011;     //93pi/512
   sin[94]  =  9'b110111010;     //94pi/512
   cos[94]  =  9'b001101011;     //94pi/512
   sin[95]  =  9'b110111010;     //95pi/512
   cos[95]  =  9'b001101010;     //95pi/512
   sin[96]  =  9'b110111001;     //96pi/512
   cos[96]  =  9'b001101010;     //96pi/512
   sin[97]  =  9'b110111000;     //97pi/512
   cos[97]  =  9'b001101001;     //97pi/512
   sin[98]  =  9'b110111000;     //98pi/512
   cos[98]  =  9'b001101001;     //98pi/512
   sin[99]  =  9'b110110111;     //99pi/512
   cos[99]  =  9'b001101001;     //99pi/512
   sin[100]  =  9'b110110110;     //100pi/512
   cos[100]  =  9'b001101000;     //100pi/512
   sin[101]  =  9'b110110110;     //101pi/512
   cos[101]  =  9'b001101000;     //101pi/512
   sin[102]  =  9'b110110101;     //102pi/512
   cos[102]  =  9'b001100111;     //102pi/512
   sin[103]  =  9'b110110100;     //103pi/512
   cos[103]  =  9'b001100111;     //103pi/512
   sin[104]  =  9'b110110100;     //104pi/512
   cos[104]  =  9'b001100110;     //104pi/512
   sin[105]  =  9'b110110011;     //105pi/512
   cos[105]  =  9'b001100110;     //105pi/512
   sin[106]  =  9'b110110010;     //106pi/512
   cos[106]  =  9'b001100101;     //106pi/512
   sin[107]  =  9'b110110010;     //107pi/512
   cos[107]  =  9'b001100101;     //107pi/512
   sin[108]  =  9'b110110001;     //108pi/512
   cos[108]  =  9'b001100100;     //108pi/512
   sin[109]  =  9'b110110001;     //109pi/512
   cos[109]  =  9'b001100100;     //109pi/512
   sin[110]  =  9'b110110000;     //110pi/512
   cos[110]  =  9'b001100011;     //110pi/512
   sin[111]  =  9'b110101111;     //111pi/512
   cos[111]  =  9'b001100011;     //111pi/512
   sin[112]  =  9'b110101111;     //112pi/512
   cos[112]  =  9'b001100010;     //112pi/512
   sin[113]  =  9'b110101110;     //113pi/512
   cos[113]  =  9'b001100010;     //113pi/512
   sin[114]  =  9'b110101110;     //114pi/512
   cos[114]  =  9'b001100001;     //114pi/512
   sin[115]  =  9'b110101101;     //115pi/512
   cos[115]  =  9'b001100001;     //115pi/512
   sin[116]  =  9'b110101100;     //116pi/512
   cos[116]  =  9'b001100000;     //116pi/512
   sin[117]  =  9'b110101100;     //117pi/512
   cos[117]  =  9'b001100000;     //117pi/512
   sin[118]  =  9'b110101011;     //118pi/512
   cos[118]  =  9'b001011111;     //118pi/512
   sin[119]  =  9'b110101011;     //119pi/512
   cos[119]  =  9'b001011111;     //119pi/512
   sin[120]  =  9'b110101010;     //120pi/512
   cos[120]  =  9'b001011110;     //120pi/512
   sin[121]  =  9'b110101001;     //121pi/512
   cos[121]  =  9'b001011110;     //121pi/512
   sin[122]  =  9'b110101001;     //122pi/512
   cos[122]  =  9'b001011101;     //122pi/512
   sin[123]  =  9'b110101000;     //123pi/512
   cos[123]  =  9'b001011101;     //123pi/512
   sin[124]  =  9'b110101000;     //124pi/512
   cos[124]  =  9'b001011100;     //124pi/512
   sin[125]  =  9'b110100111;     //125pi/512
   cos[125]  =  9'b001011100;     //125pi/512
   sin[126]  =  9'b110100111;     //126pi/512
   cos[126]  =  9'b001011011;     //126pi/512
   sin[127]  =  9'b110100110;     //127pi/512
   cos[127]  =  9'b001011011;     //127pi/512
   sin[128]  =  9'b110100101;     //128pi/512
   cos[128]  =  9'b001011010;     //128pi/512
   sin[129]  =  9'b110100101;     //129pi/512
   cos[129]  =  9'b001011001;     //129pi/512
   sin[130]  =  9'b110100100;     //130pi/512
   cos[130]  =  9'b001011001;     //130pi/512
   sin[131]  =  9'b110100100;     //131pi/512
   cos[131]  =  9'b001011000;     //131pi/512
   sin[132]  =  9'b110100011;     //132pi/512
   cos[132]  =  9'b001011000;     //132pi/512
   sin[133]  =  9'b110100011;     //133pi/512
   cos[133]  =  9'b001010111;     //133pi/512
   sin[134]  =  9'b110100010;     //134pi/512
   cos[134]  =  9'b001010111;     //134pi/512
   sin[135]  =  9'b110100010;     //135pi/512
   cos[135]  =  9'b001010110;     //135pi/512
   sin[136]  =  9'b110100001;     //136pi/512
   cos[136]  =  9'b001010101;     //136pi/512
   sin[137]  =  9'b110100001;     //137pi/512
   cos[137]  =  9'b001010101;     //137pi/512
   sin[138]  =  9'b110100000;     //138pi/512
   cos[138]  =  9'b001010100;     //138pi/512
   sin[139]  =  9'b110100000;     //139pi/512
   cos[139]  =  9'b001010100;     //139pi/512
   sin[140]  =  9'b110011111;     //140pi/512
   cos[140]  =  9'b001010011;     //140pi/512
   sin[141]  =  9'b110011111;     //141pi/512
   cos[141]  =  9'b001010011;     //141pi/512
   sin[142]  =  9'b110011110;     //142pi/512
   cos[142]  =  9'b001010010;     //142pi/512
   sin[143]  =  9'b110011110;     //143pi/512
   cos[143]  =  9'b001010001;     //143pi/512
   sin[144]  =  9'b110011101;     //144pi/512
   cos[144]  =  9'b001010001;     //144pi/512
   sin[145]  =  9'b110011101;     //145pi/512
   cos[145]  =  9'b001010000;     //145pi/512
   sin[146]  =  9'b110011100;     //146pi/512
   cos[146]  =  9'b001001111;     //146pi/512
   sin[147]  =  9'b110011100;     //147pi/512
   cos[147]  =  9'b001001111;     //147pi/512
   sin[148]  =  9'b110011011;     //148pi/512
   cos[148]  =  9'b001001110;     //148pi/512
   sin[149]  =  9'b110011011;     //149pi/512
   cos[149]  =  9'b001001110;     //149pi/512
   sin[150]  =  9'b110011010;     //150pi/512
   cos[150]  =  9'b001001101;     //150pi/512
   sin[151]  =  9'b110011010;     //151pi/512
   cos[151]  =  9'b001001100;     //151pi/512
   sin[152]  =  9'b110011001;     //152pi/512
   cos[152]  =  9'b001001100;     //152pi/512
   sin[153]  =  9'b110011001;     //153pi/512
   cos[153]  =  9'b001001011;     //153pi/512
   sin[154]  =  9'b110011000;     //154pi/512
   cos[154]  =  9'b001001010;     //154pi/512
   sin[155]  =  9'b110011000;     //155pi/512
   cos[155]  =  9'b001001010;     //155pi/512
   sin[156]  =  9'b110010111;     //156pi/512
   cos[156]  =  9'b001001001;     //156pi/512
   sin[157]  =  9'b110010111;     //157pi/512
   cos[157]  =  9'b001001001;     //157pi/512
   sin[158]  =  9'b110010110;     //158pi/512
   cos[158]  =  9'b001001000;     //158pi/512
   sin[159]  =  9'b110010110;     //159pi/512
   cos[159]  =  9'b001000111;     //159pi/512
   sin[160]  =  9'b110010110;     //160pi/512
   cos[160]  =  9'b001000111;     //160pi/512
   sin[161]  =  9'b110010101;     //161pi/512
   cos[161]  =  9'b001000110;     //161pi/512
   sin[162]  =  9'b110010101;     //162pi/512
   cos[162]  =  9'b001000101;     //162pi/512
   sin[163]  =  9'b110010100;     //163pi/512
   cos[163]  =  9'b001000101;     //163pi/512
   sin[164]  =  9'b110010100;     //164pi/512
   cos[164]  =  9'b001000100;     //164pi/512
   sin[165]  =  9'b110010011;     //165pi/512
   cos[165]  =  9'b001000011;     //165pi/512
   sin[166]  =  9'b110010011;     //166pi/512
   cos[166]  =  9'b001000011;     //166pi/512
   sin[167]  =  9'b110010011;     //167pi/512
   cos[167]  =  9'b001000010;     //167pi/512
   sin[168]  =  9'b110010010;     //168pi/512
   cos[168]  =  9'b001000001;     //168pi/512
   sin[169]  =  9'b110010010;     //169pi/512
   cos[169]  =  9'b001000001;     //169pi/512
   sin[170]  =  9'b110010001;     //170pi/512
   cos[170]  =  9'b001000000;     //170pi/512
   sin[171]  =  9'b110010001;     //171pi/512
   cos[171]  =  9'b000111111;     //171pi/512
   sin[172]  =  9'b110010001;     //172pi/512
   cos[172]  =  9'b000111111;     //172pi/512
   sin[173]  =  9'b110010000;     //173pi/512
   cos[173]  =  9'b000111110;     //173pi/512
   sin[174]  =  9'b110010000;     //174pi/512
   cos[174]  =  9'b000111101;     //174pi/512
   sin[175]  =  9'b110001111;     //175pi/512
   cos[175]  =  9'b000111101;     //175pi/512
   sin[176]  =  9'b110001111;     //176pi/512
   cos[176]  =  9'b000111100;     //176pi/512
   sin[177]  =  9'b110001111;     //177pi/512
   cos[177]  =  9'b000111011;     //177pi/512
   sin[178]  =  9'b110001110;     //178pi/512
   cos[178]  =  9'b000111010;     //178pi/512
   sin[179]  =  9'b110001110;     //179pi/512
   cos[179]  =  9'b000111010;     //179pi/512
   sin[180]  =  9'b110001110;     //180pi/512
   cos[180]  =  9'b000111001;     //180pi/512
   sin[181]  =  9'b110001101;     //181pi/512
   cos[181]  =  9'b000111000;     //181pi/512
   sin[182]  =  9'b110001101;     //182pi/512
   cos[182]  =  9'b000111000;     //182pi/512
   sin[183]  =  9'b110001101;     //183pi/512
   cos[183]  =  9'b000110111;     //183pi/512
   sin[184]  =  9'b110001100;     //184pi/512
   cos[184]  =  9'b000110110;     //184pi/512
   sin[185]  =  9'b110001100;     //185pi/512
   cos[185]  =  9'b000110110;     //185pi/512
   sin[186]  =  9'b110001100;     //186pi/512
   cos[186]  =  9'b000110101;     //186pi/512
   sin[187]  =  9'b110001011;     //187pi/512
   cos[187]  =  9'b000110100;     //187pi/512
   sin[188]  =  9'b110001011;     //188pi/512
   cos[188]  =  9'b000110011;     //188pi/512
   sin[189]  =  9'b110001011;     //189pi/512
   cos[189]  =  9'b000110011;     //189pi/512
   sin[190]  =  9'b110001010;     //190pi/512
   cos[190]  =  9'b000110010;     //190pi/512
   sin[191]  =  9'b110001010;     //191pi/512
   cos[191]  =  9'b000110001;     //191pi/512
   sin[192]  =  9'b110001010;     //192pi/512
   cos[192]  =  9'b000110000;     //192pi/512
   sin[193]  =  9'b110001001;     //193pi/512
   cos[193]  =  9'b000110000;     //193pi/512
   sin[194]  =  9'b110001001;     //194pi/512
   cos[194]  =  9'b000101111;     //194pi/512
   sin[195]  =  9'b110001001;     //195pi/512
   cos[195]  =  9'b000101110;     //195pi/512
   sin[196]  =  9'b110001001;     //196pi/512
   cos[196]  =  9'b000101110;     //196pi/512
   sin[197]  =  9'b110001000;     //197pi/512
   cos[197]  =  9'b000101101;     //197pi/512
   sin[198]  =  9'b110001000;     //198pi/512
   cos[198]  =  9'b000101100;     //198pi/512
   sin[199]  =  9'b110001000;     //199pi/512
   cos[199]  =  9'b000101011;     //199pi/512
   sin[200]  =  9'b110000111;     //200pi/512
   cos[200]  =  9'b000101011;     //200pi/512
   sin[201]  =  9'b110000111;     //201pi/512
   cos[201]  =  9'b000101010;     //201pi/512
   sin[202]  =  9'b110000111;     //202pi/512
   cos[202]  =  9'b000101001;     //202pi/512
   sin[203]  =  9'b110000111;     //203pi/512
   cos[203]  =  9'b000101000;     //203pi/512
   sin[204]  =  9'b110000110;     //204pi/512
   cos[204]  =  9'b000101000;     //204pi/512
   sin[205]  =  9'b110000110;     //205pi/512
   cos[205]  =  9'b000100111;     //205pi/512
   sin[206]  =  9'b110000110;     //206pi/512
   cos[206]  =  9'b000100110;     //206pi/512
   sin[207]  =  9'b110000110;     //207pi/512
   cos[207]  =  9'b000100101;     //207pi/512
   sin[208]  =  9'b110000110;     //208pi/512
   cos[208]  =  9'b000100101;     //208pi/512
   sin[209]  =  9'b110000101;     //209pi/512
   cos[209]  =  9'b000100100;     //209pi/512
   sin[210]  =  9'b110000101;     //210pi/512
   cos[210]  =  9'b000100011;     //210pi/512
   sin[211]  =  9'b110000101;     //211pi/512
   cos[211]  =  9'b000100010;     //211pi/512
   sin[212]  =  9'b110000101;     //212pi/512
   cos[212]  =  9'b000100010;     //212pi/512
   sin[213]  =  9'b110000100;     //213pi/512
   cos[213]  =  9'b000100001;     //213pi/512
   sin[214]  =  9'b110000100;     //214pi/512
   cos[214]  =  9'b000100000;     //214pi/512
   sin[215]  =  9'b110000100;     //215pi/512
   cos[215]  =  9'b000011111;     //215pi/512
   sin[216]  =  9'b110000100;     //216pi/512
   cos[216]  =  9'b000011111;     //216pi/512
   sin[217]  =  9'b110000100;     //217pi/512
   cos[217]  =  9'b000011110;     //217pi/512
   sin[218]  =  9'b110000011;     //218pi/512
   cos[218]  =  9'b000011101;     //218pi/512
   sin[219]  =  9'b110000011;     //219pi/512
   cos[219]  =  9'b000011100;     //219pi/512
   sin[220]  =  9'b110000011;     //220pi/512
   cos[220]  =  9'b000011100;     //220pi/512
   sin[221]  =  9'b110000011;     //221pi/512
   cos[221]  =  9'b000011011;     //221pi/512
   sin[222]  =  9'b110000011;     //222pi/512
   cos[222]  =  9'b000011010;     //222pi/512
   sin[223]  =  9'b110000011;     //223pi/512
   cos[223]  =  9'b000011001;     //223pi/512
   sin[224]  =  9'b110000010;     //224pi/512
   cos[224]  =  9'b000011000;     //224pi/512
   sin[225]  =  9'b110000010;     //225pi/512
   cos[225]  =  9'b000011000;     //225pi/512
   sin[226]  =  9'b110000010;     //226pi/512
   cos[226]  =  9'b000010111;     //226pi/512
   sin[227]  =  9'b110000010;     //227pi/512
   cos[227]  =  9'b000010110;     //227pi/512
   sin[228]  =  9'b110000010;     //228pi/512
   cos[228]  =  9'b000010101;     //228pi/512
   sin[229]  =  9'b110000010;     //229pi/512
   cos[229]  =  9'b000010101;     //229pi/512
   sin[230]  =  9'b110000010;     //230pi/512
   cos[230]  =  9'b000010100;     //230pi/512
   sin[231]  =  9'b110000010;     //231pi/512
   cos[231]  =  9'b000010011;     //231pi/512
   sin[232]  =  9'b110000001;     //232pi/512
   cos[232]  =  9'b000010010;     //232pi/512
   sin[233]  =  9'b110000001;     //233pi/512
   cos[233]  =  9'b000010010;     //233pi/512
   sin[234]  =  9'b110000001;     //234pi/512
   cos[234]  =  9'b000010001;     //234pi/512
   sin[235]  =  9'b110000001;     //235pi/512
   cos[235]  =  9'b000010000;     //235pi/512
   sin[236]  =  9'b110000001;     //236pi/512
   cos[236]  =  9'b000001111;     //236pi/512
   sin[237]  =  9'b110000001;     //237pi/512
   cos[237]  =  9'b000001110;     //237pi/512
   sin[238]  =  9'b110000001;     //238pi/512
   cos[238]  =  9'b000001110;     //238pi/512
   sin[239]  =  9'b110000001;     //239pi/512
   cos[239]  =  9'b000001101;     //239pi/512
   sin[240]  =  9'b110000001;     //240pi/512
   cos[240]  =  9'b000001100;     //240pi/512
   sin[241]  =  9'b110000001;     //241pi/512
   cos[241]  =  9'b000001011;     //241pi/512
   sin[242]  =  9'b110000000;     //242pi/512
   cos[242]  =  9'b000001010;     //242pi/512
   sin[243]  =  9'b110000000;     //243pi/512
   cos[243]  =  9'b000001010;     //243pi/512
   sin[244]  =  9'b110000000;     //244pi/512
   cos[244]  =  9'b000001001;     //244pi/512
   sin[245]  =  9'b110000000;     //245pi/512
   cos[245]  =  9'b000001000;     //245pi/512
   sin[246]  =  9'b110000000;     //246pi/512
   cos[246]  =  9'b000000111;     //246pi/512
   sin[247]  =  9'b110000000;     //247pi/512
   cos[247]  =  9'b000000111;     //247pi/512
   sin[248]  =  9'b110000000;     //248pi/512
   cos[248]  =  9'b000000110;     //248pi/512
   sin[249]  =  9'b110000000;     //249pi/512
   cos[249]  =  9'b000000101;     //249pi/512
   sin[250]  =  9'b110000000;     //250pi/512
   cos[250]  =  9'b000000100;     //250pi/512
   sin[251]  =  9'b110000000;     //251pi/512
   cos[251]  =  9'b000000011;     //251pi/512
   sin[252]  =  9'b110000000;     //252pi/512
   cos[252]  =  9'b000000011;     //252pi/512
   sin[253]  =  9'b110000000;     //253pi/512
   cos[253]  =  9'b000000010;     //253pi/512
   sin[254]  =  9'b110000000;     //254pi/512
   cos[254]  =  9'b000000001;     //254pi/512
   sin[255]  =  9'b110000000;     //255pi/512
   cos[255]  =  9'b000000000;     //255pi/512
   sin[256]  =  9'b110000000;     //256pi/512
   cos[256]  =  9'b000000000;     //256pi/512
   sin[257]  =  9'b110000000;     //257pi/512
   cos[257]  =  9'b111111111;     //257pi/512
   sin[258]  =  9'b110000000;     //258pi/512
   cos[258]  =  9'b111111110;     //258pi/512
   sin[259]  =  9'b110000000;     //259pi/512
   cos[259]  =  9'b111111110;     //259pi/512
   sin[260]  =  9'b110000000;     //260pi/512
   cos[260]  =  9'b111111101;     //260pi/512
   sin[261]  =  9'b110000000;     //261pi/512
   cos[261]  =  9'b111111100;     //261pi/512
   sin[262]  =  9'b110000000;     //262pi/512
   cos[262]  =  9'b111111011;     //262pi/512
   sin[263]  =  9'b110000000;     //263pi/512
   cos[263]  =  9'b111111011;     //263pi/512
   sin[264]  =  9'b110000000;     //264pi/512
   cos[264]  =  9'b111111010;     //264pi/512
   sin[265]  =  9'b110000000;     //265pi/512
   cos[265]  =  9'b111111001;     //265pi/512
   sin[266]  =  9'b110000000;     //266pi/512
   cos[266]  =  9'b111111000;     //266pi/512
   sin[267]  =  9'b110000000;     //267pi/512
   cos[267]  =  9'b111110111;     //267pi/512
   sin[268]  =  9'b110000000;     //268pi/512
   cos[268]  =  9'b111110111;     //268pi/512
   sin[269]  =  9'b110000000;     //269pi/512
   cos[269]  =  9'b111110110;     //269pi/512
   sin[270]  =  9'b110000000;     //270pi/512
   cos[270]  =  9'b111110101;     //270pi/512
   sin[271]  =  9'b110000001;     //271pi/512
   cos[271]  =  9'b111110100;     //271pi/512
   sin[272]  =  9'b110000001;     //272pi/512
   cos[272]  =  9'b111110011;     //272pi/512
   sin[273]  =  9'b110000001;     //273pi/512
   cos[273]  =  9'b111110011;     //273pi/512
   sin[274]  =  9'b110000001;     //274pi/512
   cos[274]  =  9'b111110010;     //274pi/512
   sin[275]  =  9'b110000001;     //275pi/512
   cos[275]  =  9'b111110001;     //275pi/512
   sin[276]  =  9'b110000001;     //276pi/512
   cos[276]  =  9'b111110000;     //276pi/512
   sin[277]  =  9'b110000001;     //277pi/512
   cos[277]  =  9'b111110000;     //277pi/512
   sin[278]  =  9'b110000001;     //278pi/512
   cos[278]  =  9'b111101111;     //278pi/512
   sin[279]  =  9'b110000001;     //279pi/512
   cos[279]  =  9'b111101110;     //279pi/512
   sin[280]  =  9'b110000001;     //280pi/512
   cos[280]  =  9'b111101101;     //280pi/512
   sin[281]  =  9'b110000010;     //281pi/512
   cos[281]  =  9'b111101100;     //281pi/512
   sin[282]  =  9'b110000010;     //282pi/512
   cos[282]  =  9'b111101100;     //282pi/512
   sin[283]  =  9'b110000010;     //283pi/512
   cos[283]  =  9'b111101011;     //283pi/512
   sin[284]  =  9'b110000010;     //284pi/512
   cos[284]  =  9'b111101010;     //284pi/512
   sin[285]  =  9'b110000010;     //285pi/512
   cos[285]  =  9'b111101001;     //285pi/512
   sin[286]  =  9'b110000010;     //286pi/512
   cos[286]  =  9'b111101001;     //286pi/512
   sin[287]  =  9'b110000010;     //287pi/512
   cos[287]  =  9'b111101000;     //287pi/512
   sin[288]  =  9'b110000010;     //288pi/512
   cos[288]  =  9'b111100111;     //288pi/512
   sin[289]  =  9'b110000011;     //289pi/512
   cos[289]  =  9'b111100110;     //289pi/512
   sin[290]  =  9'b110000011;     //290pi/512
   cos[290]  =  9'b111100101;     //290pi/512
   sin[291]  =  9'b110000011;     //291pi/512
   cos[291]  =  9'b111100101;     //291pi/512
   sin[292]  =  9'b110000011;     //292pi/512
   cos[292]  =  9'b111100100;     //292pi/512
   sin[293]  =  9'b110000011;     //293pi/512
   cos[293]  =  9'b111100011;     //293pi/512
   sin[294]  =  9'b110000011;     //294pi/512
   cos[294]  =  9'b111100010;     //294pi/512
   sin[295]  =  9'b110000100;     //295pi/512
   cos[295]  =  9'b111100010;     //295pi/512
   sin[296]  =  9'b110000100;     //296pi/512
   cos[296]  =  9'b111100001;     //296pi/512
   sin[297]  =  9'b110000100;     //297pi/512
   cos[297]  =  9'b111100000;     //297pi/512
   sin[298]  =  9'b110000100;     //298pi/512
   cos[298]  =  9'b111011111;     //298pi/512
   sin[299]  =  9'b110000100;     //299pi/512
   cos[299]  =  9'b111011111;     //299pi/512
   sin[300]  =  9'b110000101;     //300pi/512
   cos[300]  =  9'b111011110;     //300pi/512
   sin[301]  =  9'b110000101;     //301pi/512
   cos[301]  =  9'b111011101;     //301pi/512
   sin[302]  =  9'b110000101;     //302pi/512
   cos[302]  =  9'b111011100;     //302pi/512
   sin[303]  =  9'b110000101;     //303pi/512
   cos[303]  =  9'b111011100;     //303pi/512
   sin[304]  =  9'b110000110;     //304pi/512
   cos[304]  =  9'b111011011;     //304pi/512
   sin[305]  =  9'b110000110;     //305pi/512
   cos[305]  =  9'b111011010;     //305pi/512
   sin[306]  =  9'b110000110;     //306pi/512
   cos[306]  =  9'b111011001;     //306pi/512
   sin[307]  =  9'b110000110;     //307pi/512
   cos[307]  =  9'b111011001;     //307pi/512
   sin[308]  =  9'b110000110;     //308pi/512
   cos[308]  =  9'b111011000;     //308pi/512
   sin[309]  =  9'b110000111;     //309pi/512
   cos[309]  =  9'b111010111;     //309pi/512
   sin[310]  =  9'b110000111;     //310pi/512
   cos[310]  =  9'b111010110;     //310pi/512
   sin[311]  =  9'b110000111;     //311pi/512
   cos[311]  =  9'b111010110;     //311pi/512
   sin[312]  =  9'b110000111;     //312pi/512
   cos[312]  =  9'b111010101;     //312pi/512
   sin[313]  =  9'b110001000;     //313pi/512
   cos[313]  =  9'b111010100;     //313pi/512
   sin[314]  =  9'b110001000;     //314pi/512
   cos[314]  =  9'b111010011;     //314pi/512
   sin[315]  =  9'b110001000;     //315pi/512
   cos[315]  =  9'b111010011;     //315pi/512
   sin[316]  =  9'b110001001;     //316pi/512
   cos[316]  =  9'b111010010;     //316pi/512
   sin[317]  =  9'b110001001;     //317pi/512
   cos[317]  =  9'b111010001;     //317pi/512
   sin[318]  =  9'b110001001;     //318pi/512
   cos[318]  =  9'b111010000;     //318pi/512
   sin[319]  =  9'b110001001;     //319pi/512
   cos[319]  =  9'b111010000;     //319pi/512
   sin[320]  =  9'b110001010;     //320pi/512
   cos[320]  =  9'b111001111;     //320pi/512
   sin[321]  =  9'b110001010;     //321pi/512
   cos[321]  =  9'b111001110;     //321pi/512
   sin[322]  =  9'b110001010;     //322pi/512
   cos[322]  =  9'b111001110;     //322pi/512
   sin[323]  =  9'b110001011;     //323pi/512
   cos[323]  =  9'b111001101;     //323pi/512
   sin[324]  =  9'b110001011;     //324pi/512
   cos[324]  =  9'b111001100;     //324pi/512
   sin[325]  =  9'b110001011;     //325pi/512
   cos[325]  =  9'b111001011;     //325pi/512
   sin[326]  =  9'b110001100;     //326pi/512
   cos[326]  =  9'b111001011;     //326pi/512
   sin[327]  =  9'b110001100;     //327pi/512
   cos[327]  =  9'b111001010;     //327pi/512
   sin[328]  =  9'b110001100;     //328pi/512
   cos[328]  =  9'b111001001;     //328pi/512
   sin[329]  =  9'b110001101;     //329pi/512
   cos[329]  =  9'b111001001;     //329pi/512
   sin[330]  =  9'b110001101;     //330pi/512
   cos[330]  =  9'b111001000;     //330pi/512
   sin[331]  =  9'b110001101;     //331pi/512
   cos[331]  =  9'b111000111;     //331pi/512
   sin[332]  =  9'b110001110;     //332pi/512
   cos[332]  =  9'b111000110;     //332pi/512
   sin[333]  =  9'b110001110;     //333pi/512
   cos[333]  =  9'b111000110;     //333pi/512
   sin[334]  =  9'b110001110;     //334pi/512
   cos[334]  =  9'b111000101;     //334pi/512
   sin[335]  =  9'b110001111;     //335pi/512
   cos[335]  =  9'b111000100;     //335pi/512
   sin[336]  =  9'b110001111;     //336pi/512
   cos[336]  =  9'b111000100;     //336pi/512
   sin[337]  =  9'b110001111;     //337pi/512
   cos[337]  =  9'b111000011;     //337pi/512
   sin[338]  =  9'b110010000;     //338pi/512
   cos[338]  =  9'b111000010;     //338pi/512
   sin[339]  =  9'b110010000;     //339pi/512
   cos[339]  =  9'b111000010;     //339pi/512
   sin[340]  =  9'b110010001;     //340pi/512
   cos[340]  =  9'b111000001;     //340pi/512
   sin[341]  =  9'b110010001;     //341pi/512
   cos[341]  =  9'b111000000;     //341pi/512
   sin[342]  =  9'b110010001;     //342pi/512
   cos[342]  =  9'b111000000;     //342pi/512
   sin[343]  =  9'b110010010;     //343pi/512
   cos[343]  =  9'b110111111;     //343pi/512
   sin[344]  =  9'b110010010;     //344pi/512
   cos[344]  =  9'b110111110;     //344pi/512
   sin[345]  =  9'b110010011;     //345pi/512
   cos[345]  =  9'b110111110;     //345pi/512
   sin[346]  =  9'b110010011;     //346pi/512
   cos[346]  =  9'b110111101;     //346pi/512
   sin[347]  =  9'b110010011;     //347pi/512
   cos[347]  =  9'b110111100;     //347pi/512
   sin[348]  =  9'b110010100;     //348pi/512
   cos[348]  =  9'b110111100;     //348pi/512
   sin[349]  =  9'b110010100;     //349pi/512
   cos[349]  =  9'b110111011;     //349pi/512
   sin[350]  =  9'b110010101;     //350pi/512
   cos[350]  =  9'b110111010;     //350pi/512
   sin[351]  =  9'b110010101;     //351pi/512
   cos[351]  =  9'b110111010;     //351pi/512
   sin[352]  =  9'b110010110;     //352pi/512
   cos[352]  =  9'b110111001;     //352pi/512
   sin[353]  =  9'b110010110;     //353pi/512
   cos[353]  =  9'b110111000;     //353pi/512
   sin[354]  =  9'b110010110;     //354pi/512
   cos[354]  =  9'b110111000;     //354pi/512
   sin[355]  =  9'b110010111;     //355pi/512
   cos[355]  =  9'b110110111;     //355pi/512
   sin[356]  =  9'b110010111;     //356pi/512
   cos[356]  =  9'b110110110;     //356pi/512
   sin[357]  =  9'b110011000;     //357pi/512
   cos[357]  =  9'b110110110;     //357pi/512
   sin[358]  =  9'b110011000;     //358pi/512
   cos[358]  =  9'b110110101;     //358pi/512
   sin[359]  =  9'b110011001;     //359pi/512
   cos[359]  =  9'b110110100;     //359pi/512
   sin[360]  =  9'b110011001;     //360pi/512
   cos[360]  =  9'b110110100;     //360pi/512
   sin[361]  =  9'b110011010;     //361pi/512
   cos[361]  =  9'b110110011;     //361pi/512
   sin[362]  =  9'b110011010;     //362pi/512
   cos[362]  =  9'b110110010;     //362pi/512
   sin[363]  =  9'b110011011;     //363pi/512
   cos[363]  =  9'b110110010;     //363pi/512
   sin[364]  =  9'b110011011;     //364pi/512
   cos[364]  =  9'b110110001;     //364pi/512
   sin[365]  =  9'b110011100;     //365pi/512
   cos[365]  =  9'b110110001;     //365pi/512
   sin[366]  =  9'b110011100;     //366pi/512
   cos[366]  =  9'b110110000;     //366pi/512
   sin[367]  =  9'b110011101;     //367pi/512
   cos[367]  =  9'b110101111;     //367pi/512
   sin[368]  =  9'b110011101;     //368pi/512
   cos[368]  =  9'b110101111;     //368pi/512
   sin[369]  =  9'b110011110;     //369pi/512
   cos[369]  =  9'b110101110;     //369pi/512
   sin[370]  =  9'b110011110;     //370pi/512
   cos[370]  =  9'b110101110;     //370pi/512
   sin[371]  =  9'b110011111;     //371pi/512
   cos[371]  =  9'b110101101;     //371pi/512
   sin[372]  =  9'b110011111;     //372pi/512
   cos[372]  =  9'b110101100;     //372pi/512
   sin[373]  =  9'b110100000;     //373pi/512
   cos[373]  =  9'b110101100;     //373pi/512
   sin[374]  =  9'b110100000;     //374pi/512
   cos[374]  =  9'b110101011;     //374pi/512
   sin[375]  =  9'b110100001;     //375pi/512
   cos[375]  =  9'b110101011;     //375pi/512
   sin[376]  =  9'b110100001;     //376pi/512
   cos[376]  =  9'b110101010;     //376pi/512
   sin[377]  =  9'b110100010;     //377pi/512
   cos[377]  =  9'b110101001;     //377pi/512
   sin[378]  =  9'b110100010;     //378pi/512
   cos[378]  =  9'b110101001;     //378pi/512
   sin[379]  =  9'b110100011;     //379pi/512
   cos[379]  =  9'b110101000;     //379pi/512
   sin[380]  =  9'b110100011;     //380pi/512
   cos[380]  =  9'b110101000;     //380pi/512
   sin[381]  =  9'b110100100;     //381pi/512
   cos[381]  =  9'b110100111;     //381pi/512
   sin[382]  =  9'b110100100;     //382pi/512
   cos[382]  =  9'b110100111;     //382pi/512
   sin[383]  =  9'b110100101;     //383pi/512
   cos[383]  =  9'b110100110;     //383pi/512
   sin[384]  =  9'b110100101;     //384pi/512
   cos[384]  =  9'b110100101;     //384pi/512
   sin[385]  =  9'b110100110;     //385pi/512
   cos[385]  =  9'b110100101;     //385pi/512
   sin[386]  =  9'b110100111;     //386pi/512
   cos[386]  =  9'b110100100;     //386pi/512
   sin[387]  =  9'b110100111;     //387pi/512
   cos[387]  =  9'b110100100;     //387pi/512
   sin[388]  =  9'b110101000;     //388pi/512
   cos[388]  =  9'b110100011;     //388pi/512
   sin[389]  =  9'b110101000;     //389pi/512
   cos[389]  =  9'b110100011;     //389pi/512
   sin[390]  =  9'b110101001;     //390pi/512
   cos[390]  =  9'b110100010;     //390pi/512
   sin[391]  =  9'b110101001;     //391pi/512
   cos[391]  =  9'b110100010;     //391pi/512
   sin[392]  =  9'b110101010;     //392pi/512
   cos[392]  =  9'b110100001;     //392pi/512
   sin[393]  =  9'b110101011;     //393pi/512
   cos[393]  =  9'b110100001;     //393pi/512
   sin[394]  =  9'b110101011;     //394pi/512
   cos[394]  =  9'b110100000;     //394pi/512
   sin[395]  =  9'b110101100;     //395pi/512
   cos[395]  =  9'b110100000;     //395pi/512
   sin[396]  =  9'b110101100;     //396pi/512
   cos[396]  =  9'b110011111;     //396pi/512
   sin[397]  =  9'b110101101;     //397pi/512
   cos[397]  =  9'b110011111;     //397pi/512
   sin[398]  =  9'b110101110;     //398pi/512
   cos[398]  =  9'b110011110;     //398pi/512
   sin[399]  =  9'b110101110;     //399pi/512
   cos[399]  =  9'b110011110;     //399pi/512
   sin[400]  =  9'b110101111;     //400pi/512
   cos[400]  =  9'b110011101;     //400pi/512
   sin[401]  =  9'b110101111;     //401pi/512
   cos[401]  =  9'b110011101;     //401pi/512
   sin[402]  =  9'b110110000;     //402pi/512
   cos[402]  =  9'b110011100;     //402pi/512
   sin[403]  =  9'b110110001;     //403pi/512
   cos[403]  =  9'b110011100;     //403pi/512
   sin[404]  =  9'b110110001;     //404pi/512
   cos[404]  =  9'b110011011;     //404pi/512
   sin[405]  =  9'b110110010;     //405pi/512
   cos[405]  =  9'b110011011;     //405pi/512
   sin[406]  =  9'b110110010;     //406pi/512
   cos[406]  =  9'b110011010;     //406pi/512
   sin[407]  =  9'b110110011;     //407pi/512
   cos[407]  =  9'b110011010;     //407pi/512
   sin[408]  =  9'b110110100;     //408pi/512
   cos[408]  =  9'b110011001;     //408pi/512
   sin[409]  =  9'b110110100;     //409pi/512
   cos[409]  =  9'b110011001;     //409pi/512
   sin[410]  =  9'b110110101;     //410pi/512
   cos[410]  =  9'b110011000;     //410pi/512
   sin[411]  =  9'b110110110;     //411pi/512
   cos[411]  =  9'b110011000;     //411pi/512
   sin[412]  =  9'b110110110;     //412pi/512
   cos[412]  =  9'b110010111;     //412pi/512
   sin[413]  =  9'b110110111;     //413pi/512
   cos[413]  =  9'b110010111;     //413pi/512
   sin[414]  =  9'b110111000;     //414pi/512
   cos[414]  =  9'b110010110;     //414pi/512
   sin[415]  =  9'b110111000;     //415pi/512
   cos[415]  =  9'b110010110;     //415pi/512
   sin[416]  =  9'b110111001;     //416pi/512
   cos[416]  =  9'b110010110;     //416pi/512
   sin[417]  =  9'b110111010;     //417pi/512
   cos[417]  =  9'b110010101;     //417pi/512
   sin[418]  =  9'b110111010;     //418pi/512
   cos[418]  =  9'b110010101;     //418pi/512
   sin[419]  =  9'b110111011;     //419pi/512
   cos[419]  =  9'b110010100;     //419pi/512
   sin[420]  =  9'b110111100;     //420pi/512
   cos[420]  =  9'b110010100;     //420pi/512
   sin[421]  =  9'b110111100;     //421pi/512
   cos[421]  =  9'b110010011;     //421pi/512
   sin[422]  =  9'b110111101;     //422pi/512
   cos[422]  =  9'b110010011;     //422pi/512
   sin[423]  =  9'b110111110;     //423pi/512
   cos[423]  =  9'b110010011;     //423pi/512
   sin[424]  =  9'b110111110;     //424pi/512
   cos[424]  =  9'b110010010;     //424pi/512
   sin[425]  =  9'b110111111;     //425pi/512
   cos[425]  =  9'b110010010;     //425pi/512
   sin[426]  =  9'b111000000;     //426pi/512
   cos[426]  =  9'b110010001;     //426pi/512
   sin[427]  =  9'b111000000;     //427pi/512
   cos[427]  =  9'b110010001;     //427pi/512
   sin[428]  =  9'b111000001;     //428pi/512
   cos[428]  =  9'b110010001;     //428pi/512
   sin[429]  =  9'b111000010;     //429pi/512
   cos[429]  =  9'b110010000;     //429pi/512
   sin[430]  =  9'b111000010;     //430pi/512
   cos[430]  =  9'b110010000;     //430pi/512
   sin[431]  =  9'b111000011;     //431pi/512
   cos[431]  =  9'b110001111;     //431pi/512
   sin[432]  =  9'b111000100;     //432pi/512
   cos[432]  =  9'b110001111;     //432pi/512
   sin[433]  =  9'b111000100;     //433pi/512
   cos[433]  =  9'b110001111;     //433pi/512
   sin[434]  =  9'b111000101;     //434pi/512
   cos[434]  =  9'b110001110;     //434pi/512
   sin[435]  =  9'b111000110;     //435pi/512
   cos[435]  =  9'b110001110;     //435pi/512
   sin[436]  =  9'b111000110;     //436pi/512
   cos[436]  =  9'b110001110;     //436pi/512
   sin[437]  =  9'b111000111;     //437pi/512
   cos[437]  =  9'b110001101;     //437pi/512
   sin[438]  =  9'b111001000;     //438pi/512
   cos[438]  =  9'b110001101;     //438pi/512
   sin[439]  =  9'b111001001;     //439pi/512
   cos[439]  =  9'b110001101;     //439pi/512
   sin[440]  =  9'b111001001;     //440pi/512
   cos[440]  =  9'b110001100;     //440pi/512
   sin[441]  =  9'b111001010;     //441pi/512
   cos[441]  =  9'b110001100;     //441pi/512
   sin[442]  =  9'b111001011;     //442pi/512
   cos[442]  =  9'b110001100;     //442pi/512
   sin[443]  =  9'b111001011;     //443pi/512
   cos[443]  =  9'b110001011;     //443pi/512
   sin[444]  =  9'b111001100;     //444pi/512
   cos[444]  =  9'b110001011;     //444pi/512
   sin[445]  =  9'b111001101;     //445pi/512
   cos[445]  =  9'b110001011;     //445pi/512
   sin[446]  =  9'b111001110;     //446pi/512
   cos[446]  =  9'b110001010;     //446pi/512
   sin[447]  =  9'b111001110;     //447pi/512
   cos[447]  =  9'b110001010;     //447pi/512
   sin[448]  =  9'b111001111;     //448pi/512
   cos[448]  =  9'b110001010;     //448pi/512
   sin[449]  =  9'b111010000;     //449pi/512
   cos[449]  =  9'b110001001;     //449pi/512
   sin[450]  =  9'b111010000;     //450pi/512
   cos[450]  =  9'b110001001;     //450pi/512
   sin[451]  =  9'b111010001;     //451pi/512
   cos[451]  =  9'b110001001;     //451pi/512
   sin[452]  =  9'b111010010;     //452pi/512
   cos[452]  =  9'b110001001;     //452pi/512
   sin[453]  =  9'b111010011;     //453pi/512
   cos[453]  =  9'b110001000;     //453pi/512
   sin[454]  =  9'b111010011;     //454pi/512
   cos[454]  =  9'b110001000;     //454pi/512
   sin[455]  =  9'b111010100;     //455pi/512
   cos[455]  =  9'b110001000;     //455pi/512
   sin[456]  =  9'b111010101;     //456pi/512
   cos[456]  =  9'b110000111;     //456pi/512
   sin[457]  =  9'b111010110;     //457pi/512
   cos[457]  =  9'b110000111;     //457pi/512
   sin[458]  =  9'b111010110;     //458pi/512
   cos[458]  =  9'b110000111;     //458pi/512
   sin[459]  =  9'b111010111;     //459pi/512
   cos[459]  =  9'b110000111;     //459pi/512
   sin[460]  =  9'b111011000;     //460pi/512
   cos[460]  =  9'b110000110;     //460pi/512
   sin[461]  =  9'b111011001;     //461pi/512
   cos[461]  =  9'b110000110;     //461pi/512
   sin[462]  =  9'b111011001;     //462pi/512
   cos[462]  =  9'b110000110;     //462pi/512
   sin[463]  =  9'b111011010;     //463pi/512
   cos[463]  =  9'b110000110;     //463pi/512
   sin[464]  =  9'b111011011;     //464pi/512
   cos[464]  =  9'b110000110;     //464pi/512
   sin[465]  =  9'b111011100;     //465pi/512
   cos[465]  =  9'b110000101;     //465pi/512
   sin[466]  =  9'b111011100;     //466pi/512
   cos[466]  =  9'b110000101;     //466pi/512
   sin[467]  =  9'b111011101;     //467pi/512
   cos[467]  =  9'b110000101;     //467pi/512
   sin[468]  =  9'b111011110;     //468pi/512
   cos[468]  =  9'b110000101;     //468pi/512
   sin[469]  =  9'b111011111;     //469pi/512
   cos[469]  =  9'b110000100;     //469pi/512
   sin[470]  =  9'b111011111;     //470pi/512
   cos[470]  =  9'b110000100;     //470pi/512
   sin[471]  =  9'b111100000;     //471pi/512
   cos[471]  =  9'b110000100;     //471pi/512
   sin[472]  =  9'b111100001;     //472pi/512
   cos[472]  =  9'b110000100;     //472pi/512
   sin[473]  =  9'b111100010;     //473pi/512
   cos[473]  =  9'b110000100;     //473pi/512
   sin[474]  =  9'b111100010;     //474pi/512
   cos[474]  =  9'b110000011;     //474pi/512
   sin[475]  =  9'b111100011;     //475pi/512
   cos[475]  =  9'b110000011;     //475pi/512
   sin[476]  =  9'b111100100;     //476pi/512
   cos[476]  =  9'b110000011;     //476pi/512
   sin[477]  =  9'b111100101;     //477pi/512
   cos[477]  =  9'b110000011;     //477pi/512
   sin[478]  =  9'b111100101;     //478pi/512
   cos[478]  =  9'b110000011;     //478pi/512
   sin[479]  =  9'b111100110;     //479pi/512
   cos[479]  =  9'b110000011;     //479pi/512
   sin[480]  =  9'b111100111;     //480pi/512
   cos[480]  =  9'b110000010;     //480pi/512
   sin[481]  =  9'b111101000;     //481pi/512
   cos[481]  =  9'b110000010;     //481pi/512
   sin[482]  =  9'b111101001;     //482pi/512
   cos[482]  =  9'b110000010;     //482pi/512
   sin[483]  =  9'b111101001;     //483pi/512
   cos[483]  =  9'b110000010;     //483pi/512
   sin[484]  =  9'b111101010;     //484pi/512
   cos[484]  =  9'b110000010;     //484pi/512
   sin[485]  =  9'b111101011;     //485pi/512
   cos[485]  =  9'b110000010;     //485pi/512
   sin[486]  =  9'b111101100;     //486pi/512
   cos[486]  =  9'b110000010;     //486pi/512
   sin[487]  =  9'b111101100;     //487pi/512
   cos[487]  =  9'b110000010;     //487pi/512
   sin[488]  =  9'b111101101;     //488pi/512
   cos[488]  =  9'b110000001;     //488pi/512
   sin[489]  =  9'b111101110;     //489pi/512
   cos[489]  =  9'b110000001;     //489pi/512
   sin[490]  =  9'b111101111;     //490pi/512
   cos[490]  =  9'b110000001;     //490pi/512
   sin[491]  =  9'b111110000;     //491pi/512
   cos[491]  =  9'b110000001;     //491pi/512
   sin[492]  =  9'b111110000;     //492pi/512
   cos[492]  =  9'b110000001;     //492pi/512
   sin[493]  =  9'b111110001;     //493pi/512
   cos[493]  =  9'b110000001;     //493pi/512
   sin[494]  =  9'b111110010;     //494pi/512
   cos[494]  =  9'b110000001;     //494pi/512
   sin[495]  =  9'b111110011;     //495pi/512
   cos[495]  =  9'b110000001;     //495pi/512
   sin[496]  =  9'b111110011;     //496pi/512
   cos[496]  =  9'b110000001;     //496pi/512
   sin[497]  =  9'b111110100;     //497pi/512
   cos[497]  =  9'b110000001;     //497pi/512
   sin[498]  =  9'b111110101;     //498pi/512
   cos[498]  =  9'b110000000;     //498pi/512
   sin[499]  =  9'b111110110;     //499pi/512
   cos[499]  =  9'b110000000;     //499pi/512
   sin[500]  =  9'b111110111;     //500pi/512
   cos[500]  =  9'b110000000;     //500pi/512
   sin[501]  =  9'b111110111;     //501pi/512
   cos[501]  =  9'b110000000;     //501pi/512
   sin[502]  =  9'b111111000;     //502pi/512
   cos[502]  =  9'b110000000;     //502pi/512
   sin[503]  =  9'b111111001;     //503pi/512
   cos[503]  =  9'b110000000;     //503pi/512
   sin[504]  =  9'b111111010;     //504pi/512
   cos[504]  =  9'b110000000;     //504pi/512
   sin[505]  =  9'b111111011;     //505pi/512
   cos[505]  =  9'b110000000;     //505pi/512
   sin[506]  =  9'b111111011;     //506pi/512
   cos[506]  =  9'b110000000;     //506pi/512
   sin[507]  =  9'b111111100;     //507pi/512
   cos[507]  =  9'b110000000;     //507pi/512
   sin[508]  =  9'b111111101;     //508pi/512
   cos[508]  =  9'b110000000;     //508pi/512
   sin[509]  =  9'b111111110;     //509pi/512
   cos[509]  =  9'b110000000;     //509pi/512
   sin[510]  =  9'b111111110;     //510pi/512
   cos[510]  =  9'b110000000;     //510pi/512
   sin[511]  =  9'b111111111;     //511pi/512
   cos[511]  =  9'b110000000;     //511pi/512
end
endmodule