module  M_TWIDLE_11_B_0_5_v  #(parameter SIZE = 10, word_length_tw = 11) (
    input            clk,
    input            en_rd,
    input   [10:0]   rd_ptr_angle,
    input            en_modf,
    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );
reg signed [word_length_tw-1:0]  cos    [511:0];
reg signed [word_length_tw-1:0]  sin    [511:0];
reg signed [word_length_tw-1:0]  m_cos  [511:0];
reg signed [word_length_tw-1:0]  m_sin  [511:0];
reg signed [word_length_tw-1:0]  cos_temp;
reg signed [word_length_tw-1:0]  sin_temp;
reg signed [word_length_tw-1:0]  m_cos_temp;
reg signed [word_length_tw-1:0]  m_sin_temp;
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & ~ en_modf) begin
                  cos_temp           <= cos   [rd_ptr_angle];
                  sin_temp           <= sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & en_modf) begin
                  m_cos_temp           <= m_cos   [rd_ptr_angle];
                  m_sin_temp           <= m_sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(*) begin 
             if (en_modf) begin
                  cos_data           <= m_cos_temp;
                  sin_data           <= m_sin_temp;
             end else begin
                  cos_data           <= cos_temp;
                  sin_data           <= sin_temp;
             end 
        end
initial begin
   sin[0]  =  11'b00000000000;     //0pi/512
   cos[0]  =  11'b01000000000;     //0pi/512
   sin[1]  =  11'b11111111101;     //1pi/512
   cos[1]  =  11'b00111111111;     //1pi/512
   sin[2]  =  11'b11111111010;     //2pi/512
   cos[2]  =  11'b00111111111;     //2pi/512
   sin[3]  =  11'b11111110111;     //3pi/512
   cos[3]  =  11'b00111111111;     //3pi/512
   sin[4]  =  11'b11111110011;     //4pi/512
   cos[4]  =  11'b00111111111;     //4pi/512
   sin[5]  =  11'b11111110000;     //5pi/512
   cos[5]  =  11'b00111111111;     //5pi/512
   sin[6]  =  11'b11111101101;     //6pi/512
   cos[6]  =  11'b00111111111;     //6pi/512
   sin[7]  =  11'b11111101010;     //7pi/512
   cos[7]  =  11'b00111111111;     //7pi/512
   sin[8]  =  11'b11111100111;     //8pi/512
   cos[8]  =  11'b00111111111;     //8pi/512
   sin[9]  =  11'b11111100100;     //9pi/512
   cos[9]  =  11'b00111111111;     //9pi/512
   sin[10]  =  11'b11111100001;     //10pi/512
   cos[10]  =  11'b00111111111;     //10pi/512
   sin[11]  =  11'b11111011101;     //11pi/512
   cos[11]  =  11'b00111111110;     //11pi/512
   sin[12]  =  11'b11111011010;     //12pi/512
   cos[12]  =  11'b00111111110;     //12pi/512
   sin[13]  =  11'b11111010111;     //13pi/512
   cos[13]  =  11'b00111111110;     //13pi/512
   sin[14]  =  11'b11111010100;     //14pi/512
   cos[14]  =  11'b00111111110;     //14pi/512
   sin[15]  =  11'b11111010001;     //15pi/512
   cos[15]  =  11'b00111111101;     //15pi/512
   sin[16]  =  11'b11111001110;     //16pi/512
   cos[16]  =  11'b00111111101;     //16pi/512
   sin[17]  =  11'b11111001011;     //17pi/512
   cos[17]  =  11'b00111111101;     //17pi/512
   sin[18]  =  11'b11111001000;     //18pi/512
   cos[18]  =  11'b00111111100;     //18pi/512
   sin[19]  =  11'b11111000100;     //19pi/512
   cos[19]  =  11'b00111111100;     //19pi/512
   sin[20]  =  11'b11111000001;     //20pi/512
   cos[20]  =  11'b00111111100;     //20pi/512
   sin[21]  =  11'b11110111110;     //21pi/512
   cos[21]  =  11'b00111111011;     //21pi/512
   sin[22]  =  11'b11110111011;     //22pi/512
   cos[22]  =  11'b00111111011;     //22pi/512
   sin[23]  =  11'b11110111000;     //23pi/512
   cos[23]  =  11'b00111111010;     //23pi/512
   sin[24]  =  11'b11110110101;     //24pi/512
   cos[24]  =  11'b00111111010;     //24pi/512
   sin[25]  =  11'b11110110010;     //25pi/512
   cos[25]  =  11'b00111111001;     //25pi/512
   sin[26]  =  11'b11110101111;     //26pi/512
   cos[26]  =  11'b00111111001;     //26pi/512
   sin[27]  =  11'b11110101100;     //27pi/512
   cos[27]  =  11'b00111111000;     //27pi/512
   sin[28]  =  11'b11110101000;     //28pi/512
   cos[28]  =  11'b00111111000;     //28pi/512
   sin[29]  =  11'b11110100101;     //29pi/512
   cos[29]  =  11'b00111110111;     //29pi/512
   sin[30]  =  11'b11110100010;     //30pi/512
   cos[30]  =  11'b00111110111;     //30pi/512
   sin[31]  =  11'b11110011111;     //31pi/512
   cos[31]  =  11'b00111110110;     //31pi/512
   sin[32]  =  11'b11110011100;     //32pi/512
   cos[32]  =  11'b00111110110;     //32pi/512
   sin[33]  =  11'b11110011001;     //33pi/512
   cos[33]  =  11'b00111110101;     //33pi/512
   sin[34]  =  11'b11110010110;     //34pi/512
   cos[34]  =  11'b00111110100;     //34pi/512
   sin[35]  =  11'b11110010011;     //35pi/512
   cos[35]  =  11'b00111110100;     //35pi/512
   sin[36]  =  11'b11110010000;     //36pi/512
   cos[36]  =  11'b00111110011;     //36pi/512
   sin[37]  =  11'b11110001101;     //37pi/512
   cos[37]  =  11'b00111110010;     //37pi/512
   sin[38]  =  11'b11110001010;     //38pi/512
   cos[38]  =  11'b00111110010;     //38pi/512
   sin[39]  =  11'b11110000111;     //39pi/512
   cos[39]  =  11'b00111110001;     //39pi/512
   sin[40]  =  11'b11110000100;     //40pi/512
   cos[40]  =  11'b00111110000;     //40pi/512
   sin[41]  =  11'b11110000001;     //41pi/512
   cos[41]  =  11'b00111101111;     //41pi/512
   sin[42]  =  11'b11101111110;     //42pi/512
   cos[42]  =  11'b00111101111;     //42pi/512
   sin[43]  =  11'b11101111010;     //43pi/512
   cos[43]  =  11'b00111101110;     //43pi/512
   sin[44]  =  11'b11101110111;     //44pi/512
   cos[44]  =  11'b00111101101;     //44pi/512
   sin[45]  =  11'b11101110100;     //45pi/512
   cos[45]  =  11'b00111101100;     //45pi/512
   sin[46]  =  11'b11101110001;     //46pi/512
   cos[46]  =  11'b00111101011;     //46pi/512
   sin[47]  =  11'b11101101110;     //47pi/512
   cos[47]  =  11'b00111101010;     //47pi/512
   sin[48]  =  11'b11101101011;     //48pi/512
   cos[48]  =  11'b00111101001;     //48pi/512
   sin[49]  =  11'b11101101000;     //49pi/512
   cos[49]  =  11'b00111101001;     //49pi/512
   sin[50]  =  11'b11101100101;     //50pi/512
   cos[50]  =  11'b00111101000;     //50pi/512
   sin[51]  =  11'b11101100010;     //51pi/512
   cos[51]  =  11'b00111100111;     //51pi/512
   sin[52]  =  11'b11101011111;     //52pi/512
   cos[52]  =  11'b00111100110;     //52pi/512
   sin[53]  =  11'b11101011100;     //53pi/512
   cos[53]  =  11'b00111100101;     //53pi/512
   sin[54]  =  11'b11101011001;     //54pi/512
   cos[54]  =  11'b00111100100;     //54pi/512
   sin[55]  =  11'b11101010110;     //55pi/512
   cos[55]  =  11'b00111100011;     //55pi/512
   sin[56]  =  11'b11101010100;     //56pi/512
   cos[56]  =  11'b00111100010;     //56pi/512
   sin[57]  =  11'b11101010001;     //57pi/512
   cos[57]  =  11'b00111100001;     //57pi/512
   sin[58]  =  11'b11101001110;     //58pi/512
   cos[58]  =  11'b00111011111;     //58pi/512
   sin[59]  =  11'b11101001011;     //59pi/512
   cos[59]  =  11'b00111011110;     //59pi/512
   sin[60]  =  11'b11101001000;     //60pi/512
   cos[60]  =  11'b00111011101;     //60pi/512
   sin[61]  =  11'b11101000101;     //61pi/512
   cos[61]  =  11'b00111011100;     //61pi/512
   sin[62]  =  11'b11101000010;     //62pi/512
   cos[62]  =  11'b00111011011;     //62pi/512
   sin[63]  =  11'b11100111111;     //63pi/512
   cos[63]  =  11'b00111011010;     //63pi/512
   sin[64]  =  11'b11100111100;     //64pi/512
   cos[64]  =  11'b00111011001;     //64pi/512
   sin[65]  =  11'b11100111001;     //65pi/512
   cos[65]  =  11'b00111010111;     //65pi/512
   sin[66]  =  11'b11100110110;     //66pi/512
   cos[66]  =  11'b00111010110;     //66pi/512
   sin[67]  =  11'b11100110011;     //67pi/512
   cos[67]  =  11'b00111010101;     //67pi/512
   sin[68]  =  11'b11100110001;     //68pi/512
   cos[68]  =  11'b00111010100;     //68pi/512
   sin[69]  =  11'b11100101110;     //69pi/512
   cos[69]  =  11'b00111010010;     //69pi/512
   sin[70]  =  11'b11100101011;     //70pi/512
   cos[70]  =  11'b00111010001;     //70pi/512
   sin[71]  =  11'b11100101000;     //71pi/512
   cos[71]  =  11'b00111010000;     //71pi/512
   sin[72]  =  11'b11100100101;     //72pi/512
   cos[72]  =  11'b00111001110;     //72pi/512
   sin[73]  =  11'b11100100010;     //73pi/512
   cos[73]  =  11'b00111001101;     //73pi/512
   sin[74]  =  11'b11100011111;     //74pi/512
   cos[74]  =  11'b00111001100;     //74pi/512
   sin[75]  =  11'b11100011101;     //75pi/512
   cos[75]  =  11'b00111001010;     //75pi/512
   sin[76]  =  11'b11100011010;     //76pi/512
   cos[76]  =  11'b00111001001;     //76pi/512
   sin[77]  =  11'b11100010111;     //77pi/512
   cos[77]  =  11'b00111000111;     //77pi/512
   sin[78]  =  11'b11100010100;     //78pi/512
   cos[78]  =  11'b00111000110;     //78pi/512
   sin[79]  =  11'b11100010001;     //79pi/512
   cos[79]  =  11'b00111000101;     //79pi/512
   sin[80]  =  11'b11100001111;     //80pi/512
   cos[80]  =  11'b00111000011;     //80pi/512
   sin[81]  =  11'b11100001100;     //81pi/512
   cos[81]  =  11'b00111000010;     //81pi/512
   sin[82]  =  11'b11100001001;     //82pi/512
   cos[82]  =  11'b00111000000;     //82pi/512
   sin[83]  =  11'b11100000110;     //83pi/512
   cos[83]  =  11'b00110111111;     //83pi/512
   sin[84]  =  11'b11100000100;     //84pi/512
   cos[84]  =  11'b00110111101;     //84pi/512
   sin[85]  =  11'b11100000001;     //85pi/512
   cos[85]  =  11'b00110111011;     //85pi/512
   sin[86]  =  11'b11011111110;     //86pi/512
   cos[86]  =  11'b00110111010;     //86pi/512
   sin[87]  =  11'b11011111011;     //87pi/512
   cos[87]  =  11'b00110111000;     //87pi/512
   sin[88]  =  11'b11011111001;     //88pi/512
   cos[88]  =  11'b00110110111;     //88pi/512
   sin[89]  =  11'b11011110110;     //89pi/512
   cos[89]  =  11'b00110110101;     //89pi/512
   sin[90]  =  11'b11011110011;     //90pi/512
   cos[90]  =  11'b00110110011;     //90pi/512
   sin[91]  =  11'b11011110001;     //91pi/512
   cos[91]  =  11'b00110110010;     //91pi/512
   sin[92]  =  11'b11011101110;     //92pi/512
   cos[92]  =  11'b00110110000;     //92pi/512
   sin[93]  =  11'b11011101011;     //93pi/512
   cos[93]  =  11'b00110101110;     //93pi/512
   sin[94]  =  11'b11011101001;     //94pi/512
   cos[94]  =  11'b00110101101;     //94pi/512
   sin[95]  =  11'b11011100110;     //95pi/512
   cos[95]  =  11'b00110101011;     //95pi/512
   sin[96]  =  11'b11011100100;     //96pi/512
   cos[96]  =  11'b00110101001;     //96pi/512
   sin[97]  =  11'b11011100001;     //97pi/512
   cos[97]  =  11'b00110100111;     //97pi/512
   sin[98]  =  11'b11011011110;     //98pi/512
   cos[98]  =  11'b00110100110;     //98pi/512
   sin[99]  =  11'b11011011100;     //99pi/512
   cos[99]  =  11'b00110100100;     //99pi/512
   sin[100]  =  11'b11011011001;     //100pi/512
   cos[100]  =  11'b00110100010;     //100pi/512
   sin[101]  =  11'b11011010111;     //101pi/512
   cos[101]  =  11'b00110100000;     //101pi/512
   sin[102]  =  11'b11011010100;     //102pi/512
   cos[102]  =  11'b00110011110;     //102pi/512
   sin[103]  =  11'b11011010010;     //103pi/512
   cos[103]  =  11'b00110011101;     //103pi/512
   sin[104]  =  11'b11011001111;     //104pi/512
   cos[104]  =  11'b00110011011;     //104pi/512
   sin[105]  =  11'b11011001100;     //105pi/512
   cos[105]  =  11'b00110011001;     //105pi/512
   sin[106]  =  11'b11011001010;     //106pi/512
   cos[106]  =  11'b00110010111;     //106pi/512
   sin[107]  =  11'b11011000111;     //107pi/512
   cos[107]  =  11'b00110010101;     //107pi/512
   sin[108]  =  11'b11011000101;     //108pi/512
   cos[108]  =  11'b00110010011;     //108pi/512
   sin[109]  =  11'b11011000011;     //109pi/512
   cos[109]  =  11'b00110010001;     //109pi/512
   sin[110]  =  11'b11011000000;     //110pi/512
   cos[110]  =  11'b00110001111;     //110pi/512
   sin[111]  =  11'b11010111110;     //111pi/512
   cos[111]  =  11'b00110001101;     //111pi/512
   sin[112]  =  11'b11010111011;     //112pi/512
   cos[112]  =  11'b00110001011;     //112pi/512
   sin[113]  =  11'b11010111001;     //113pi/512
   cos[113]  =  11'b00110001001;     //113pi/512
   sin[114]  =  11'b11010110110;     //114pi/512
   cos[114]  =  11'b00110000111;     //114pi/512
   sin[115]  =  11'b11010110100;     //115pi/512
   cos[115]  =  11'b00110000101;     //115pi/512
   sin[116]  =  11'b11010110010;     //116pi/512
   cos[116]  =  11'b00110000011;     //116pi/512
   sin[117]  =  11'b11010101111;     //117pi/512
   cos[117]  =  11'b00110000001;     //117pi/512
   sin[118]  =  11'b11010101101;     //118pi/512
   cos[118]  =  11'b00101111111;     //118pi/512
   sin[119]  =  11'b11010101010;     //119pi/512
   cos[119]  =  11'b00101111101;     //119pi/512
   sin[120]  =  11'b11010101000;     //120pi/512
   cos[120]  =  11'b00101111011;     //120pi/512
   sin[121]  =  11'b11010100110;     //121pi/512
   cos[121]  =  11'b00101111001;     //121pi/512
   sin[122]  =  11'b11010100100;     //122pi/512
   cos[122]  =  11'b00101110111;     //122pi/512
   sin[123]  =  11'b11010100001;     //123pi/512
   cos[123]  =  11'b00101110100;     //123pi/512
   sin[124]  =  11'b11010011111;     //124pi/512
   cos[124]  =  11'b00101110010;     //124pi/512
   sin[125]  =  11'b11010011101;     //125pi/512
   cos[125]  =  11'b00101110000;     //125pi/512
   sin[126]  =  11'b11010011010;     //126pi/512
   cos[126]  =  11'b00101101110;     //126pi/512
   sin[127]  =  11'b11010011000;     //127pi/512
   cos[127]  =  11'b00101101100;     //127pi/512
   sin[128]  =  11'b11010010110;     //128pi/512
   cos[128]  =  11'b00101101010;     //128pi/512
   sin[129]  =  11'b11010010100;     //129pi/512
   cos[129]  =  11'b00101100111;     //129pi/512
   sin[130]  =  11'b11010010010;     //130pi/512
   cos[130]  =  11'b00101100101;     //130pi/512
   sin[131]  =  11'b11010001111;     //131pi/512
   cos[131]  =  11'b00101100011;     //131pi/512
   sin[132]  =  11'b11010001101;     //132pi/512
   cos[132]  =  11'b00101100001;     //132pi/512
   sin[133]  =  11'b11010001011;     //133pi/512
   cos[133]  =  11'b00101011110;     //133pi/512
   sin[134]  =  11'b11010001001;     //134pi/512
   cos[134]  =  11'b00101011100;     //134pi/512
   sin[135]  =  11'b11010000111;     //135pi/512
   cos[135]  =  11'b00101011010;     //135pi/512
   sin[136]  =  11'b11010000101;     //136pi/512
   cos[136]  =  11'b00101010111;     //136pi/512
   sin[137]  =  11'b11010000011;     //137pi/512
   cos[137]  =  11'b00101010101;     //137pi/512
   sin[138]  =  11'b11010000000;     //138pi/512
   cos[138]  =  11'b00101010011;     //138pi/512
   sin[139]  =  11'b11001111110;     //139pi/512
   cos[139]  =  11'b00101010000;     //139pi/512
   sin[140]  =  11'b11001111100;     //140pi/512
   cos[140]  =  11'b00101001110;     //140pi/512
   sin[141]  =  11'b11001111010;     //141pi/512
   cos[141]  =  11'b00101001100;     //141pi/512
   sin[142]  =  11'b11001111000;     //142pi/512
   cos[142]  =  11'b00101001001;     //142pi/512
   sin[143]  =  11'b11001110110;     //143pi/512
   cos[143]  =  11'b00101000111;     //143pi/512
   sin[144]  =  11'b11001110100;     //144pi/512
   cos[144]  =  11'b00101000100;     //144pi/512
   sin[145]  =  11'b11001110010;     //145pi/512
   cos[145]  =  11'b00101000010;     //145pi/512
   sin[146]  =  11'b11001110000;     //146pi/512
   cos[146]  =  11'b00100111111;     //146pi/512
   sin[147]  =  11'b11001101110;     //147pi/512
   cos[147]  =  11'b00100111101;     //147pi/512
   sin[148]  =  11'b11001101100;     //148pi/512
   cos[148]  =  11'b00100111010;     //148pi/512
   sin[149]  =  11'b11001101010;     //149pi/512
   cos[149]  =  11'b00100111000;     //149pi/512
   sin[150]  =  11'b11001101001;     //150pi/512
   cos[150]  =  11'b00100110110;     //150pi/512
   sin[151]  =  11'b11001100111;     //151pi/512
   cos[151]  =  11'b00100110011;     //151pi/512
   sin[152]  =  11'b11001100101;     //152pi/512
   cos[152]  =  11'b00100110000;     //152pi/512
   sin[153]  =  11'b11001100011;     //153pi/512
   cos[153]  =  11'b00100101110;     //153pi/512
   sin[154]  =  11'b11001100001;     //154pi/512
   cos[154]  =  11'b00100101011;     //154pi/512
   sin[155]  =  11'b11001011111;     //155pi/512
   cos[155]  =  11'b00100101001;     //155pi/512
   sin[156]  =  11'b11001011101;     //156pi/512
   cos[156]  =  11'b00100100110;     //156pi/512
   sin[157]  =  11'b11001011100;     //157pi/512
   cos[157]  =  11'b00100100100;     //157pi/512
   sin[158]  =  11'b11001011010;     //158pi/512
   cos[158]  =  11'b00100100001;     //158pi/512
   sin[159]  =  11'b11001011000;     //159pi/512
   cos[159]  =  11'b00100011111;     //159pi/512
   sin[160]  =  11'b11001010110;     //160pi/512
   cos[160]  =  11'b00100011100;     //160pi/512
   sin[161]  =  11'b11001010101;     //161pi/512
   cos[161]  =  11'b00100011001;     //161pi/512
   sin[162]  =  11'b11001010011;     //162pi/512
   cos[162]  =  11'b00100010111;     //162pi/512
   sin[163]  =  11'b11001010001;     //163pi/512
   cos[163]  =  11'b00100010100;     //163pi/512
   sin[164]  =  11'b11001001111;     //164pi/512
   cos[164]  =  11'b00100010001;     //164pi/512
   sin[165]  =  11'b11001001110;     //165pi/512
   cos[165]  =  11'b00100001111;     //165pi/512
   sin[166]  =  11'b11001001100;     //166pi/512
   cos[166]  =  11'b00100001100;     //166pi/512
   sin[167]  =  11'b11001001010;     //167pi/512
   cos[167]  =  11'b00100001001;     //167pi/512
   sin[168]  =  11'b11001001001;     //168pi/512
   cos[168]  =  11'b00100000111;     //168pi/512
   sin[169]  =  11'b11001000111;     //169pi/512
   cos[169]  =  11'b00100000100;     //169pi/512
   sin[170]  =  11'b11001000110;     //170pi/512
   cos[170]  =  11'b00100000001;     //170pi/512
   sin[171]  =  11'b11001000100;     //171pi/512
   cos[171]  =  11'b00011111111;     //171pi/512
   sin[172]  =  11'b11001000011;     //172pi/512
   cos[172]  =  11'b00011111100;     //172pi/512
   sin[173]  =  11'b11001000001;     //173pi/512
   cos[173]  =  11'b00011111001;     //173pi/512
   sin[174]  =  11'b11000111111;     //174pi/512
   cos[174]  =  11'b00011110110;     //174pi/512
   sin[175]  =  11'b11000111110;     //175pi/512
   cos[175]  =  11'b00011110100;     //175pi/512
   sin[176]  =  11'b11000111100;     //176pi/512
   cos[176]  =  11'b00011110001;     //176pi/512
   sin[177]  =  11'b11000111011;     //177pi/512
   cos[177]  =  11'b00011101110;     //177pi/512
   sin[178]  =  11'b11000111010;     //178pi/512
   cos[178]  =  11'b00011101011;     //178pi/512
   sin[179]  =  11'b11000111000;     //179pi/512
   cos[179]  =  11'b00011101001;     //179pi/512
   sin[180]  =  11'b11000110111;     //180pi/512
   cos[180]  =  11'b00011100110;     //180pi/512
   sin[181]  =  11'b11000110101;     //181pi/512
   cos[181]  =  11'b00011100011;     //181pi/512
   sin[182]  =  11'b11000110100;     //182pi/512
   cos[182]  =  11'b00011100000;     //182pi/512
   sin[183]  =  11'b11000110011;     //183pi/512
   cos[183]  =  11'b00011011101;     //183pi/512
   sin[184]  =  11'b11000110001;     //184pi/512
   cos[184]  =  11'b00011011010;     //184pi/512
   sin[185]  =  11'b11000110000;     //185pi/512
   cos[185]  =  11'b00011011000;     //185pi/512
   sin[186]  =  11'b11000101111;     //186pi/512
   cos[186]  =  11'b00011010101;     //186pi/512
   sin[187]  =  11'b11000101101;     //187pi/512
   cos[187]  =  11'b00011010010;     //187pi/512
   sin[188]  =  11'b11000101100;     //188pi/512
   cos[188]  =  11'b00011001111;     //188pi/512
   sin[189]  =  11'b11000101011;     //189pi/512
   cos[189]  =  11'b00011001100;     //189pi/512
   sin[190]  =  11'b11000101001;     //190pi/512
   cos[190]  =  11'b00011001001;     //190pi/512
   sin[191]  =  11'b11000101000;     //191pi/512
   cos[191]  =  11'b00011000110;     //191pi/512
   sin[192]  =  11'b11000100111;     //192pi/512
   cos[192]  =  11'b00011000011;     //192pi/512
   sin[193]  =  11'b11000100110;     //193pi/512
   cos[193]  =  11'b00011000001;     //193pi/512
   sin[194]  =  11'b11000100101;     //194pi/512
   cos[194]  =  11'b00010111110;     //194pi/512
   sin[195]  =  11'b11000100011;     //195pi/512
   cos[195]  =  11'b00010111011;     //195pi/512
   sin[196]  =  11'b11000100010;     //196pi/512
   cos[196]  =  11'b00010111000;     //196pi/512
   sin[197]  =  11'b11000100001;     //197pi/512
   cos[197]  =  11'b00010110101;     //197pi/512
   sin[198]  =  11'b11000100000;     //198pi/512
   cos[198]  =  11'b00010110010;     //198pi/512
   sin[199]  =  11'b11000011111;     //199pi/512
   cos[199]  =  11'b00010101111;     //199pi/512
   sin[200]  =  11'b11000011110;     //200pi/512
   cos[200]  =  11'b00010101100;     //200pi/512
   sin[201]  =  11'b11000011101;     //201pi/512
   cos[201]  =  11'b00010101001;     //201pi/512
   sin[202]  =  11'b11000011100;     //202pi/512
   cos[202]  =  11'b00010100110;     //202pi/512
   sin[203]  =  11'b11000011011;     //203pi/512
   cos[203]  =  11'b00010100011;     //203pi/512
   sin[204]  =  11'b11000011010;     //204pi/512
   cos[204]  =  11'b00010100000;     //204pi/512
   sin[205]  =  11'b11000011001;     //205pi/512
   cos[205]  =  11'b00010011101;     //205pi/512
   sin[206]  =  11'b11000011000;     //206pi/512
   cos[206]  =  11'b00010011010;     //206pi/512
   sin[207]  =  11'b11000010111;     //207pi/512
   cos[207]  =  11'b00010010111;     //207pi/512
   sin[208]  =  11'b11000010110;     //208pi/512
   cos[208]  =  11'b00010010100;     //208pi/512
   sin[209]  =  11'b11000010101;     //209pi/512
   cos[209]  =  11'b00010010001;     //209pi/512
   sin[210]  =  11'b11000010100;     //210pi/512
   cos[210]  =  11'b00010001110;     //210pi/512
   sin[211]  =  11'b11000010011;     //211pi/512
   cos[211]  =  11'b00010001011;     //211pi/512
   sin[212]  =  11'b11000010011;     //212pi/512
   cos[212]  =  11'b00010001000;     //212pi/512
   sin[213]  =  11'b11000010010;     //213pi/512
   cos[213]  =  11'b00010000101;     //213pi/512
   sin[214]  =  11'b11000010001;     //214pi/512
   cos[214]  =  11'b00010000010;     //214pi/512
   sin[215]  =  11'b11000010000;     //215pi/512
   cos[215]  =  11'b00001111111;     //215pi/512
   sin[216]  =  11'b11000001111;     //216pi/512
   cos[216]  =  11'b00001111100;     //216pi/512
   sin[217]  =  11'b11000001111;     //217pi/512
   cos[217]  =  11'b00001111001;     //217pi/512
   sin[218]  =  11'b11000001110;     //218pi/512
   cos[218]  =  11'b00001110110;     //218pi/512
   sin[219]  =  11'b11000001101;     //219pi/512
   cos[219]  =  11'b00001110011;     //219pi/512
   sin[220]  =  11'b11000001100;     //220pi/512
   cos[220]  =  11'b00001110000;     //220pi/512
   sin[221]  =  11'b11000001100;     //221pi/512
   cos[221]  =  11'b00001101101;     //221pi/512
   sin[222]  =  11'b11000001011;     //222pi/512
   cos[222]  =  11'b00001101010;     //222pi/512
   sin[223]  =  11'b11000001010;     //223pi/512
   cos[223]  =  11'b00001100110;     //223pi/512
   sin[224]  =  11'b11000001010;     //224pi/512
   cos[224]  =  11'b00001100011;     //224pi/512
   sin[225]  =  11'b11000001001;     //225pi/512
   cos[225]  =  11'b00001100000;     //225pi/512
   sin[226]  =  11'b11000001001;     //226pi/512
   cos[226]  =  11'b00001011101;     //226pi/512
   sin[227]  =  11'b11000001000;     //227pi/512
   cos[227]  =  11'b00001011010;     //227pi/512
   sin[228]  =  11'b11000001000;     //228pi/512
   cos[228]  =  11'b00001010111;     //228pi/512
   sin[229]  =  11'b11000000111;     //229pi/512
   cos[229]  =  11'b00001010100;     //229pi/512
   sin[230]  =  11'b11000000111;     //230pi/512
   cos[230]  =  11'b00001010001;     //230pi/512
   sin[231]  =  11'b11000000110;     //231pi/512
   cos[231]  =  11'b00001001110;     //231pi/512
   sin[232]  =  11'b11000000110;     //232pi/512
   cos[232]  =  11'b00001001011;     //232pi/512
   sin[233]  =  11'b11000000101;     //233pi/512
   cos[233]  =  11'b00001001000;     //233pi/512
   sin[234]  =  11'b11000000101;     //234pi/512
   cos[234]  =  11'b00001000100;     //234pi/512
   sin[235]  =  11'b11000000100;     //235pi/512
   cos[235]  =  11'b00001000001;     //235pi/512
   sin[236]  =  11'b11000000100;     //236pi/512
   cos[236]  =  11'b00000111110;     //236pi/512
   sin[237]  =  11'b11000000011;     //237pi/512
   cos[237]  =  11'b00000111011;     //237pi/512
   sin[238]  =  11'b11000000011;     //238pi/512
   cos[238]  =  11'b00000111000;     //238pi/512
   sin[239]  =  11'b11000000011;     //239pi/512
   cos[239]  =  11'b00000110101;     //239pi/512
   sin[240]  =  11'b11000000010;     //240pi/512
   cos[240]  =  11'b00000110010;     //240pi/512
   sin[241]  =  11'b11000000010;     //241pi/512
   cos[241]  =  11'b00000101111;     //241pi/512
   sin[242]  =  11'b11000000010;     //242pi/512
   cos[242]  =  11'b00000101011;     //242pi/512
   sin[243]  =  11'b11000000010;     //243pi/512
   cos[243]  =  11'b00000101000;     //243pi/512
   sin[244]  =  11'b11000000001;     //244pi/512
   cos[244]  =  11'b00000100101;     //244pi/512
   sin[245]  =  11'b11000000001;     //245pi/512
   cos[245]  =  11'b00000100010;     //245pi/512
   sin[246]  =  11'b11000000001;     //246pi/512
   cos[246]  =  11'b00000011111;     //246pi/512
   sin[247]  =  11'b11000000001;     //247pi/512
   cos[247]  =  11'b00000011100;     //247pi/512
   sin[248]  =  11'b11000000001;     //248pi/512
   cos[248]  =  11'b00000011001;     //248pi/512
   sin[249]  =  11'b11000000000;     //249pi/512
   cos[249]  =  11'b00000010101;     //249pi/512
   sin[250]  =  11'b11000000000;     //250pi/512
   cos[250]  =  11'b00000010010;     //250pi/512
   sin[251]  =  11'b11000000000;     //251pi/512
   cos[251]  =  11'b00000001111;     //251pi/512
   sin[252]  =  11'b11000000000;     //252pi/512
   cos[252]  =  11'b00000001100;     //252pi/512
   sin[253]  =  11'b11000000000;     //253pi/512
   cos[253]  =  11'b00000001001;     //253pi/512
   sin[254]  =  11'b11000000000;     //254pi/512
   cos[254]  =  11'b00000000110;     //254pi/512
   sin[255]  =  11'b11000000000;     //255pi/512
   cos[255]  =  11'b00000000011;     //255pi/512
   sin[256]  =  11'b11000000000;     //256pi/512
   cos[256]  =  11'b00000000000;     //256pi/512
   sin[257]  =  11'b11000000000;     //257pi/512
   cos[257]  =  11'b11111111101;     //257pi/512
   sin[258]  =  11'b11000000000;     //258pi/512
   cos[258]  =  11'b11111111010;     //258pi/512
   sin[259]  =  11'b11000000000;     //259pi/512
   cos[259]  =  11'b11111110111;     //259pi/512
   sin[260]  =  11'b11000000000;     //260pi/512
   cos[260]  =  11'b11111110011;     //260pi/512
   sin[261]  =  11'b11000000000;     //261pi/512
   cos[261]  =  11'b11111110000;     //261pi/512
   sin[262]  =  11'b11000000000;     //262pi/512
   cos[262]  =  11'b11111101101;     //262pi/512
   sin[263]  =  11'b11000000000;     //263pi/512
   cos[263]  =  11'b11111101010;     //263pi/512
   sin[264]  =  11'b11000000001;     //264pi/512
   cos[264]  =  11'b11111100111;     //264pi/512
   sin[265]  =  11'b11000000001;     //265pi/512
   cos[265]  =  11'b11111100100;     //265pi/512
   sin[266]  =  11'b11000000001;     //266pi/512
   cos[266]  =  11'b11111100001;     //266pi/512
   sin[267]  =  11'b11000000001;     //267pi/512
   cos[267]  =  11'b11111011101;     //267pi/512
   sin[268]  =  11'b11000000001;     //268pi/512
   cos[268]  =  11'b11111011010;     //268pi/512
   sin[269]  =  11'b11000000010;     //269pi/512
   cos[269]  =  11'b11111010111;     //269pi/512
   sin[270]  =  11'b11000000010;     //270pi/512
   cos[270]  =  11'b11111010100;     //270pi/512
   sin[271]  =  11'b11000000010;     //271pi/512
   cos[271]  =  11'b11111010001;     //271pi/512
   sin[272]  =  11'b11000000010;     //272pi/512
   cos[272]  =  11'b11111001110;     //272pi/512
   sin[273]  =  11'b11000000011;     //273pi/512
   cos[273]  =  11'b11111001011;     //273pi/512
   sin[274]  =  11'b11000000011;     //274pi/512
   cos[274]  =  11'b11111001000;     //274pi/512
   sin[275]  =  11'b11000000011;     //275pi/512
   cos[275]  =  11'b11111000100;     //275pi/512
   sin[276]  =  11'b11000000100;     //276pi/512
   cos[276]  =  11'b11111000001;     //276pi/512
   sin[277]  =  11'b11000000100;     //277pi/512
   cos[277]  =  11'b11110111110;     //277pi/512
   sin[278]  =  11'b11000000101;     //278pi/512
   cos[278]  =  11'b11110111011;     //278pi/512
   sin[279]  =  11'b11000000101;     //279pi/512
   cos[279]  =  11'b11110111000;     //279pi/512
   sin[280]  =  11'b11000000110;     //280pi/512
   cos[280]  =  11'b11110110101;     //280pi/512
   sin[281]  =  11'b11000000110;     //281pi/512
   cos[281]  =  11'b11110110010;     //281pi/512
   sin[282]  =  11'b11000000111;     //282pi/512
   cos[282]  =  11'b11110101111;     //282pi/512
   sin[283]  =  11'b11000000111;     //283pi/512
   cos[283]  =  11'b11110101100;     //283pi/512
   sin[284]  =  11'b11000001000;     //284pi/512
   cos[284]  =  11'b11110101000;     //284pi/512
   sin[285]  =  11'b11000001000;     //285pi/512
   cos[285]  =  11'b11110100101;     //285pi/512
   sin[286]  =  11'b11000001001;     //286pi/512
   cos[286]  =  11'b11110100010;     //286pi/512
   sin[287]  =  11'b11000001001;     //287pi/512
   cos[287]  =  11'b11110011111;     //287pi/512
   sin[288]  =  11'b11000001010;     //288pi/512
   cos[288]  =  11'b11110011100;     //288pi/512
   sin[289]  =  11'b11000001010;     //289pi/512
   cos[289]  =  11'b11110011001;     //289pi/512
   sin[290]  =  11'b11000001011;     //290pi/512
   cos[290]  =  11'b11110010110;     //290pi/512
   sin[291]  =  11'b11000001100;     //291pi/512
   cos[291]  =  11'b11110010011;     //291pi/512
   sin[292]  =  11'b11000001100;     //292pi/512
   cos[292]  =  11'b11110010000;     //292pi/512
   sin[293]  =  11'b11000001101;     //293pi/512
   cos[293]  =  11'b11110001101;     //293pi/512
   sin[294]  =  11'b11000001110;     //294pi/512
   cos[294]  =  11'b11110001010;     //294pi/512
   sin[295]  =  11'b11000001111;     //295pi/512
   cos[295]  =  11'b11110000111;     //295pi/512
   sin[296]  =  11'b11000001111;     //296pi/512
   cos[296]  =  11'b11110000100;     //296pi/512
   sin[297]  =  11'b11000010000;     //297pi/512
   cos[297]  =  11'b11110000001;     //297pi/512
   sin[298]  =  11'b11000010001;     //298pi/512
   cos[298]  =  11'b11101111110;     //298pi/512
   sin[299]  =  11'b11000010010;     //299pi/512
   cos[299]  =  11'b11101111010;     //299pi/512
   sin[300]  =  11'b11000010011;     //300pi/512
   cos[300]  =  11'b11101110111;     //300pi/512
   sin[301]  =  11'b11000010011;     //301pi/512
   cos[301]  =  11'b11101110100;     //301pi/512
   sin[302]  =  11'b11000010100;     //302pi/512
   cos[302]  =  11'b11101110001;     //302pi/512
   sin[303]  =  11'b11000010101;     //303pi/512
   cos[303]  =  11'b11101101110;     //303pi/512
   sin[304]  =  11'b11000010110;     //304pi/512
   cos[304]  =  11'b11101101011;     //304pi/512
   sin[305]  =  11'b11000010111;     //305pi/512
   cos[305]  =  11'b11101101000;     //305pi/512
   sin[306]  =  11'b11000011000;     //306pi/512
   cos[306]  =  11'b11101100101;     //306pi/512
   sin[307]  =  11'b11000011001;     //307pi/512
   cos[307]  =  11'b11101100010;     //307pi/512
   sin[308]  =  11'b11000011010;     //308pi/512
   cos[308]  =  11'b11101011111;     //308pi/512
   sin[309]  =  11'b11000011011;     //309pi/512
   cos[309]  =  11'b11101011100;     //309pi/512
   sin[310]  =  11'b11000011100;     //310pi/512
   cos[310]  =  11'b11101011001;     //310pi/512
   sin[311]  =  11'b11000011101;     //311pi/512
   cos[311]  =  11'b11101010110;     //311pi/512
   sin[312]  =  11'b11000011110;     //312pi/512
   cos[312]  =  11'b11101010100;     //312pi/512
   sin[313]  =  11'b11000011111;     //313pi/512
   cos[313]  =  11'b11101010001;     //313pi/512
   sin[314]  =  11'b11000100000;     //314pi/512
   cos[314]  =  11'b11101001110;     //314pi/512
   sin[315]  =  11'b11000100001;     //315pi/512
   cos[315]  =  11'b11101001011;     //315pi/512
   sin[316]  =  11'b11000100010;     //316pi/512
   cos[316]  =  11'b11101001000;     //316pi/512
   sin[317]  =  11'b11000100011;     //317pi/512
   cos[317]  =  11'b11101000101;     //317pi/512
   sin[318]  =  11'b11000100101;     //318pi/512
   cos[318]  =  11'b11101000010;     //318pi/512
   sin[319]  =  11'b11000100110;     //319pi/512
   cos[319]  =  11'b11100111111;     //319pi/512
   sin[320]  =  11'b11000100111;     //320pi/512
   cos[320]  =  11'b11100111100;     //320pi/512
   sin[321]  =  11'b11000101000;     //321pi/512
   cos[321]  =  11'b11100111001;     //321pi/512
   sin[322]  =  11'b11000101001;     //322pi/512
   cos[322]  =  11'b11100110110;     //322pi/512
   sin[323]  =  11'b11000101011;     //323pi/512
   cos[323]  =  11'b11100110011;     //323pi/512
   sin[324]  =  11'b11000101100;     //324pi/512
   cos[324]  =  11'b11100110001;     //324pi/512
   sin[325]  =  11'b11000101101;     //325pi/512
   cos[325]  =  11'b11100101110;     //325pi/512
   sin[326]  =  11'b11000101111;     //326pi/512
   cos[326]  =  11'b11100101011;     //326pi/512
   sin[327]  =  11'b11000110000;     //327pi/512
   cos[327]  =  11'b11100101000;     //327pi/512
   sin[328]  =  11'b11000110001;     //328pi/512
   cos[328]  =  11'b11100100101;     //328pi/512
   sin[329]  =  11'b11000110011;     //329pi/512
   cos[329]  =  11'b11100100010;     //329pi/512
   sin[330]  =  11'b11000110100;     //330pi/512
   cos[330]  =  11'b11100011111;     //330pi/512
   sin[331]  =  11'b11000110101;     //331pi/512
   cos[331]  =  11'b11100011101;     //331pi/512
   sin[332]  =  11'b11000110111;     //332pi/512
   cos[332]  =  11'b11100011010;     //332pi/512
   sin[333]  =  11'b11000111000;     //333pi/512
   cos[333]  =  11'b11100010111;     //333pi/512
   sin[334]  =  11'b11000111010;     //334pi/512
   cos[334]  =  11'b11100010100;     //334pi/512
   sin[335]  =  11'b11000111011;     //335pi/512
   cos[335]  =  11'b11100010001;     //335pi/512
   sin[336]  =  11'b11000111100;     //336pi/512
   cos[336]  =  11'b11100001111;     //336pi/512
   sin[337]  =  11'b11000111110;     //337pi/512
   cos[337]  =  11'b11100001100;     //337pi/512
   sin[338]  =  11'b11000111111;     //338pi/512
   cos[338]  =  11'b11100001001;     //338pi/512
   sin[339]  =  11'b11001000001;     //339pi/512
   cos[339]  =  11'b11100000110;     //339pi/512
   sin[340]  =  11'b11001000011;     //340pi/512
   cos[340]  =  11'b11100000100;     //340pi/512
   sin[341]  =  11'b11001000100;     //341pi/512
   cos[341]  =  11'b11100000001;     //341pi/512
   sin[342]  =  11'b11001000110;     //342pi/512
   cos[342]  =  11'b11011111110;     //342pi/512
   sin[343]  =  11'b11001000111;     //343pi/512
   cos[343]  =  11'b11011111011;     //343pi/512
   sin[344]  =  11'b11001001001;     //344pi/512
   cos[344]  =  11'b11011111001;     //344pi/512
   sin[345]  =  11'b11001001010;     //345pi/512
   cos[345]  =  11'b11011110110;     //345pi/512
   sin[346]  =  11'b11001001100;     //346pi/512
   cos[346]  =  11'b11011110011;     //346pi/512
   sin[347]  =  11'b11001001110;     //347pi/512
   cos[347]  =  11'b11011110001;     //347pi/512
   sin[348]  =  11'b11001001111;     //348pi/512
   cos[348]  =  11'b11011101110;     //348pi/512
   sin[349]  =  11'b11001010001;     //349pi/512
   cos[349]  =  11'b11011101011;     //349pi/512
   sin[350]  =  11'b11001010011;     //350pi/512
   cos[350]  =  11'b11011101001;     //350pi/512
   sin[351]  =  11'b11001010101;     //351pi/512
   cos[351]  =  11'b11011100110;     //351pi/512
   sin[352]  =  11'b11001010110;     //352pi/512
   cos[352]  =  11'b11011100100;     //352pi/512
   sin[353]  =  11'b11001011000;     //353pi/512
   cos[353]  =  11'b11011100001;     //353pi/512
   sin[354]  =  11'b11001011010;     //354pi/512
   cos[354]  =  11'b11011011110;     //354pi/512
   sin[355]  =  11'b11001011100;     //355pi/512
   cos[355]  =  11'b11011011100;     //355pi/512
   sin[356]  =  11'b11001011101;     //356pi/512
   cos[356]  =  11'b11011011001;     //356pi/512
   sin[357]  =  11'b11001011111;     //357pi/512
   cos[357]  =  11'b11011010111;     //357pi/512
   sin[358]  =  11'b11001100001;     //358pi/512
   cos[358]  =  11'b11011010100;     //358pi/512
   sin[359]  =  11'b11001100011;     //359pi/512
   cos[359]  =  11'b11011010010;     //359pi/512
   sin[360]  =  11'b11001100101;     //360pi/512
   cos[360]  =  11'b11011001111;     //360pi/512
   sin[361]  =  11'b11001100111;     //361pi/512
   cos[361]  =  11'b11011001100;     //361pi/512
   sin[362]  =  11'b11001101001;     //362pi/512
   cos[362]  =  11'b11011001010;     //362pi/512
   sin[363]  =  11'b11001101010;     //363pi/512
   cos[363]  =  11'b11011000111;     //363pi/512
   sin[364]  =  11'b11001101100;     //364pi/512
   cos[364]  =  11'b11011000101;     //364pi/512
   sin[365]  =  11'b11001101110;     //365pi/512
   cos[365]  =  11'b11011000011;     //365pi/512
   sin[366]  =  11'b11001110000;     //366pi/512
   cos[366]  =  11'b11011000000;     //366pi/512
   sin[367]  =  11'b11001110010;     //367pi/512
   cos[367]  =  11'b11010111110;     //367pi/512
   sin[368]  =  11'b11001110100;     //368pi/512
   cos[368]  =  11'b11010111011;     //368pi/512
   sin[369]  =  11'b11001110110;     //369pi/512
   cos[369]  =  11'b11010111001;     //369pi/512
   sin[370]  =  11'b11001111000;     //370pi/512
   cos[370]  =  11'b11010110110;     //370pi/512
   sin[371]  =  11'b11001111010;     //371pi/512
   cos[371]  =  11'b11010110100;     //371pi/512
   sin[372]  =  11'b11001111100;     //372pi/512
   cos[372]  =  11'b11010110010;     //372pi/512
   sin[373]  =  11'b11001111110;     //373pi/512
   cos[373]  =  11'b11010101111;     //373pi/512
   sin[374]  =  11'b11010000000;     //374pi/512
   cos[374]  =  11'b11010101101;     //374pi/512
   sin[375]  =  11'b11010000011;     //375pi/512
   cos[375]  =  11'b11010101010;     //375pi/512
   sin[376]  =  11'b11010000101;     //376pi/512
   cos[376]  =  11'b11010101000;     //376pi/512
   sin[377]  =  11'b11010000111;     //377pi/512
   cos[377]  =  11'b11010100110;     //377pi/512
   sin[378]  =  11'b11010001001;     //378pi/512
   cos[378]  =  11'b11010100100;     //378pi/512
   sin[379]  =  11'b11010001011;     //379pi/512
   cos[379]  =  11'b11010100001;     //379pi/512
   sin[380]  =  11'b11010001101;     //380pi/512
   cos[380]  =  11'b11010011111;     //380pi/512
   sin[381]  =  11'b11010001111;     //381pi/512
   cos[381]  =  11'b11010011101;     //381pi/512
   sin[382]  =  11'b11010010010;     //382pi/512
   cos[382]  =  11'b11010011010;     //382pi/512
   sin[383]  =  11'b11010010100;     //383pi/512
   cos[383]  =  11'b11010011000;     //383pi/512
   sin[384]  =  11'b11010010110;     //384pi/512
   cos[384]  =  11'b11010010110;     //384pi/512
   sin[385]  =  11'b11010011000;     //385pi/512
   cos[385]  =  11'b11010010100;     //385pi/512
   sin[386]  =  11'b11010011010;     //386pi/512
   cos[386]  =  11'b11010010010;     //386pi/512
   sin[387]  =  11'b11010011101;     //387pi/512
   cos[387]  =  11'b11010001111;     //387pi/512
   sin[388]  =  11'b11010011111;     //388pi/512
   cos[388]  =  11'b11010001101;     //388pi/512
   sin[389]  =  11'b11010100001;     //389pi/512
   cos[389]  =  11'b11010001011;     //389pi/512
   sin[390]  =  11'b11010100100;     //390pi/512
   cos[390]  =  11'b11010001001;     //390pi/512
   sin[391]  =  11'b11010100110;     //391pi/512
   cos[391]  =  11'b11010000111;     //391pi/512
   sin[392]  =  11'b11010101000;     //392pi/512
   cos[392]  =  11'b11010000101;     //392pi/512
   sin[393]  =  11'b11010101010;     //393pi/512
   cos[393]  =  11'b11010000011;     //393pi/512
   sin[394]  =  11'b11010101101;     //394pi/512
   cos[394]  =  11'b11010000000;     //394pi/512
   sin[395]  =  11'b11010101111;     //395pi/512
   cos[395]  =  11'b11001111110;     //395pi/512
   sin[396]  =  11'b11010110010;     //396pi/512
   cos[396]  =  11'b11001111100;     //396pi/512
   sin[397]  =  11'b11010110100;     //397pi/512
   cos[397]  =  11'b11001111010;     //397pi/512
   sin[398]  =  11'b11010110110;     //398pi/512
   cos[398]  =  11'b11001111000;     //398pi/512
   sin[399]  =  11'b11010111001;     //399pi/512
   cos[399]  =  11'b11001110110;     //399pi/512
   sin[400]  =  11'b11010111011;     //400pi/512
   cos[400]  =  11'b11001110100;     //400pi/512
   sin[401]  =  11'b11010111110;     //401pi/512
   cos[401]  =  11'b11001110010;     //401pi/512
   sin[402]  =  11'b11011000000;     //402pi/512
   cos[402]  =  11'b11001110000;     //402pi/512
   sin[403]  =  11'b11011000011;     //403pi/512
   cos[403]  =  11'b11001101110;     //403pi/512
   sin[404]  =  11'b11011000101;     //404pi/512
   cos[404]  =  11'b11001101100;     //404pi/512
   sin[405]  =  11'b11011000111;     //405pi/512
   cos[405]  =  11'b11001101010;     //405pi/512
   sin[406]  =  11'b11011001010;     //406pi/512
   cos[406]  =  11'b11001101001;     //406pi/512
   sin[407]  =  11'b11011001100;     //407pi/512
   cos[407]  =  11'b11001100111;     //407pi/512
   sin[408]  =  11'b11011001111;     //408pi/512
   cos[408]  =  11'b11001100101;     //408pi/512
   sin[409]  =  11'b11011010010;     //409pi/512
   cos[409]  =  11'b11001100011;     //409pi/512
   sin[410]  =  11'b11011010100;     //410pi/512
   cos[410]  =  11'b11001100001;     //410pi/512
   sin[411]  =  11'b11011010111;     //411pi/512
   cos[411]  =  11'b11001011111;     //411pi/512
   sin[412]  =  11'b11011011001;     //412pi/512
   cos[412]  =  11'b11001011101;     //412pi/512
   sin[413]  =  11'b11011011100;     //413pi/512
   cos[413]  =  11'b11001011100;     //413pi/512
   sin[414]  =  11'b11011011110;     //414pi/512
   cos[414]  =  11'b11001011010;     //414pi/512
   sin[415]  =  11'b11011100001;     //415pi/512
   cos[415]  =  11'b11001011000;     //415pi/512
   sin[416]  =  11'b11011100100;     //416pi/512
   cos[416]  =  11'b11001010110;     //416pi/512
   sin[417]  =  11'b11011100110;     //417pi/512
   cos[417]  =  11'b11001010101;     //417pi/512
   sin[418]  =  11'b11011101001;     //418pi/512
   cos[418]  =  11'b11001010011;     //418pi/512
   sin[419]  =  11'b11011101011;     //419pi/512
   cos[419]  =  11'b11001010001;     //419pi/512
   sin[420]  =  11'b11011101110;     //420pi/512
   cos[420]  =  11'b11001001111;     //420pi/512
   sin[421]  =  11'b11011110001;     //421pi/512
   cos[421]  =  11'b11001001110;     //421pi/512
   sin[422]  =  11'b11011110011;     //422pi/512
   cos[422]  =  11'b11001001100;     //422pi/512
   sin[423]  =  11'b11011110110;     //423pi/512
   cos[423]  =  11'b11001001010;     //423pi/512
   sin[424]  =  11'b11011111001;     //424pi/512
   cos[424]  =  11'b11001001001;     //424pi/512
   sin[425]  =  11'b11011111011;     //425pi/512
   cos[425]  =  11'b11001000111;     //425pi/512
   sin[426]  =  11'b11011111110;     //426pi/512
   cos[426]  =  11'b11001000110;     //426pi/512
   sin[427]  =  11'b11100000001;     //427pi/512
   cos[427]  =  11'b11001000100;     //427pi/512
   sin[428]  =  11'b11100000100;     //428pi/512
   cos[428]  =  11'b11001000011;     //428pi/512
   sin[429]  =  11'b11100000110;     //429pi/512
   cos[429]  =  11'b11001000001;     //429pi/512
   sin[430]  =  11'b11100001001;     //430pi/512
   cos[430]  =  11'b11000111111;     //430pi/512
   sin[431]  =  11'b11100001100;     //431pi/512
   cos[431]  =  11'b11000111110;     //431pi/512
   sin[432]  =  11'b11100001111;     //432pi/512
   cos[432]  =  11'b11000111100;     //432pi/512
   sin[433]  =  11'b11100010001;     //433pi/512
   cos[433]  =  11'b11000111011;     //433pi/512
   sin[434]  =  11'b11100010100;     //434pi/512
   cos[434]  =  11'b11000111010;     //434pi/512
   sin[435]  =  11'b11100010111;     //435pi/512
   cos[435]  =  11'b11000111000;     //435pi/512
   sin[436]  =  11'b11100011010;     //436pi/512
   cos[436]  =  11'b11000110111;     //436pi/512
   sin[437]  =  11'b11100011101;     //437pi/512
   cos[437]  =  11'b11000110101;     //437pi/512
   sin[438]  =  11'b11100011111;     //438pi/512
   cos[438]  =  11'b11000110100;     //438pi/512
   sin[439]  =  11'b11100100010;     //439pi/512
   cos[439]  =  11'b11000110011;     //439pi/512
   sin[440]  =  11'b11100100101;     //440pi/512
   cos[440]  =  11'b11000110001;     //440pi/512
   sin[441]  =  11'b11100101000;     //441pi/512
   cos[441]  =  11'b11000110000;     //441pi/512
   sin[442]  =  11'b11100101011;     //442pi/512
   cos[442]  =  11'b11000101111;     //442pi/512
   sin[443]  =  11'b11100101110;     //443pi/512
   cos[443]  =  11'b11000101101;     //443pi/512
   sin[444]  =  11'b11100110001;     //444pi/512
   cos[444]  =  11'b11000101100;     //444pi/512
   sin[445]  =  11'b11100110011;     //445pi/512
   cos[445]  =  11'b11000101011;     //445pi/512
   sin[446]  =  11'b11100110110;     //446pi/512
   cos[446]  =  11'b11000101001;     //446pi/512
   sin[447]  =  11'b11100111001;     //447pi/512
   cos[447]  =  11'b11000101000;     //447pi/512
   sin[448]  =  11'b11100111100;     //448pi/512
   cos[448]  =  11'b11000100111;     //448pi/512
   sin[449]  =  11'b11100111111;     //449pi/512
   cos[449]  =  11'b11000100110;     //449pi/512
   sin[450]  =  11'b11101000010;     //450pi/512
   cos[450]  =  11'b11000100101;     //450pi/512
   sin[451]  =  11'b11101000101;     //451pi/512
   cos[451]  =  11'b11000100011;     //451pi/512
   sin[452]  =  11'b11101001000;     //452pi/512
   cos[452]  =  11'b11000100010;     //452pi/512
   sin[453]  =  11'b11101001011;     //453pi/512
   cos[453]  =  11'b11000100001;     //453pi/512
   sin[454]  =  11'b11101001110;     //454pi/512
   cos[454]  =  11'b11000100000;     //454pi/512
   sin[455]  =  11'b11101010001;     //455pi/512
   cos[455]  =  11'b11000011111;     //455pi/512
   sin[456]  =  11'b11101010100;     //456pi/512
   cos[456]  =  11'b11000011110;     //456pi/512
   sin[457]  =  11'b11101010110;     //457pi/512
   cos[457]  =  11'b11000011101;     //457pi/512
   sin[458]  =  11'b11101011001;     //458pi/512
   cos[458]  =  11'b11000011100;     //458pi/512
   sin[459]  =  11'b11101011100;     //459pi/512
   cos[459]  =  11'b11000011011;     //459pi/512
   sin[460]  =  11'b11101011111;     //460pi/512
   cos[460]  =  11'b11000011010;     //460pi/512
   sin[461]  =  11'b11101100010;     //461pi/512
   cos[461]  =  11'b11000011001;     //461pi/512
   sin[462]  =  11'b11101100101;     //462pi/512
   cos[462]  =  11'b11000011000;     //462pi/512
   sin[463]  =  11'b11101101000;     //463pi/512
   cos[463]  =  11'b11000010111;     //463pi/512
   sin[464]  =  11'b11101101011;     //464pi/512
   cos[464]  =  11'b11000010110;     //464pi/512
   sin[465]  =  11'b11101101110;     //465pi/512
   cos[465]  =  11'b11000010101;     //465pi/512
   sin[466]  =  11'b11101110001;     //466pi/512
   cos[466]  =  11'b11000010100;     //466pi/512
   sin[467]  =  11'b11101110100;     //467pi/512
   cos[467]  =  11'b11000010011;     //467pi/512
   sin[468]  =  11'b11101110111;     //468pi/512
   cos[468]  =  11'b11000010011;     //468pi/512
   sin[469]  =  11'b11101111010;     //469pi/512
   cos[469]  =  11'b11000010010;     //469pi/512
   sin[470]  =  11'b11101111110;     //470pi/512
   cos[470]  =  11'b11000010001;     //470pi/512
   sin[471]  =  11'b11110000001;     //471pi/512
   cos[471]  =  11'b11000010000;     //471pi/512
   sin[472]  =  11'b11110000100;     //472pi/512
   cos[472]  =  11'b11000001111;     //472pi/512
   sin[473]  =  11'b11110000111;     //473pi/512
   cos[473]  =  11'b11000001111;     //473pi/512
   sin[474]  =  11'b11110001010;     //474pi/512
   cos[474]  =  11'b11000001110;     //474pi/512
   sin[475]  =  11'b11110001101;     //475pi/512
   cos[475]  =  11'b11000001101;     //475pi/512
   sin[476]  =  11'b11110010000;     //476pi/512
   cos[476]  =  11'b11000001100;     //476pi/512
   sin[477]  =  11'b11110010011;     //477pi/512
   cos[477]  =  11'b11000001100;     //477pi/512
   sin[478]  =  11'b11110010110;     //478pi/512
   cos[478]  =  11'b11000001011;     //478pi/512
   sin[479]  =  11'b11110011001;     //479pi/512
   cos[479]  =  11'b11000001010;     //479pi/512
   sin[480]  =  11'b11110011100;     //480pi/512
   cos[480]  =  11'b11000001010;     //480pi/512
   sin[481]  =  11'b11110011111;     //481pi/512
   cos[481]  =  11'b11000001001;     //481pi/512
   sin[482]  =  11'b11110100010;     //482pi/512
   cos[482]  =  11'b11000001001;     //482pi/512
   sin[483]  =  11'b11110100101;     //483pi/512
   cos[483]  =  11'b11000001000;     //483pi/512
   sin[484]  =  11'b11110101000;     //484pi/512
   cos[484]  =  11'b11000001000;     //484pi/512
   sin[485]  =  11'b11110101100;     //485pi/512
   cos[485]  =  11'b11000000111;     //485pi/512
   sin[486]  =  11'b11110101111;     //486pi/512
   cos[486]  =  11'b11000000111;     //486pi/512
   sin[487]  =  11'b11110110010;     //487pi/512
   cos[487]  =  11'b11000000110;     //487pi/512
   sin[488]  =  11'b11110110101;     //488pi/512
   cos[488]  =  11'b11000000110;     //488pi/512
   sin[489]  =  11'b11110111000;     //489pi/512
   cos[489]  =  11'b11000000101;     //489pi/512
   sin[490]  =  11'b11110111011;     //490pi/512
   cos[490]  =  11'b11000000101;     //490pi/512
   sin[491]  =  11'b11110111110;     //491pi/512
   cos[491]  =  11'b11000000100;     //491pi/512
   sin[492]  =  11'b11111000001;     //492pi/512
   cos[492]  =  11'b11000000100;     //492pi/512
   sin[493]  =  11'b11111000100;     //493pi/512
   cos[493]  =  11'b11000000011;     //493pi/512
   sin[494]  =  11'b11111001000;     //494pi/512
   cos[494]  =  11'b11000000011;     //494pi/512
   sin[495]  =  11'b11111001011;     //495pi/512
   cos[495]  =  11'b11000000011;     //495pi/512
   sin[496]  =  11'b11111001110;     //496pi/512
   cos[496]  =  11'b11000000010;     //496pi/512
   sin[497]  =  11'b11111010001;     //497pi/512
   cos[497]  =  11'b11000000010;     //497pi/512
   sin[498]  =  11'b11111010100;     //498pi/512
   cos[498]  =  11'b11000000010;     //498pi/512
   sin[499]  =  11'b11111010111;     //499pi/512
   cos[499]  =  11'b11000000010;     //499pi/512
   sin[500]  =  11'b11111011010;     //500pi/512
   cos[500]  =  11'b11000000001;     //500pi/512
   sin[501]  =  11'b11111011101;     //501pi/512
   cos[501]  =  11'b11000000001;     //501pi/512
   sin[502]  =  11'b11111100001;     //502pi/512
   cos[502]  =  11'b11000000001;     //502pi/512
   sin[503]  =  11'b11111100100;     //503pi/512
   cos[503]  =  11'b11000000001;     //503pi/512
   sin[504]  =  11'b11111100111;     //504pi/512
   cos[504]  =  11'b11000000001;     //504pi/512
   sin[505]  =  11'b11111101010;     //505pi/512
   cos[505]  =  11'b11000000000;     //505pi/512
   sin[506]  =  11'b11111101101;     //506pi/512
   cos[506]  =  11'b11000000000;     //506pi/512
   sin[507]  =  11'b11111110000;     //507pi/512
   cos[507]  =  11'b11000000000;     //507pi/512
   sin[508]  =  11'b11111110011;     //508pi/512
   cos[508]  =  11'b11000000000;     //508pi/512
   sin[509]  =  11'b11111110111;     //509pi/512
   cos[509]  =  11'b11000000000;     //509pi/512
   sin[510]  =  11'b11111111010;     //510pi/512
   cos[510]  =  11'b11000000000;     //510pi/512
   sin[511]  =  11'b11111111101;     //511pi/512
   cos[511]  =  11'b11000000000;     //511pi/512
   m_sin[0]  =  11'b00000000000;     //0pi/512
   m_cos[0]  =  11'b01000000000;     //0pi/512
   m_sin[1]  =  11'b11111111101;     //1pi/512
   m_cos[1]  =  11'b00111111111;     //1pi/512
   m_sin[2]  =  11'b11111111010;     //2pi/512
   m_cos[2]  =  11'b00111111111;     //2pi/512
   m_sin[3]  =  11'b11111110111;     //3pi/512
   m_cos[3]  =  11'b00111111111;     //3pi/512
   m_sin[4]  =  11'b11111110100;     //4pi/512
   m_cos[4]  =  11'b00111111111;     //4pi/512
   m_sin[5]  =  11'b11111110001;     //5pi/512
   m_cos[5]  =  11'b00111111111;     //5pi/512
   m_sin[6]  =  11'b11111101110;     //6pi/512
   m_cos[6]  =  11'b00111111111;     //6pi/512
   m_sin[7]  =  11'b11111101011;     //7pi/512
   m_cos[7]  =  11'b00111111111;     //7pi/512
   m_sin[8]  =  11'b11111101000;     //8pi/512
   m_cos[8]  =  11'b00111111111;     //8pi/512
   m_sin[9]  =  11'b11111100101;     //9pi/512
   m_cos[9]  =  11'b00111111111;     //9pi/512
   m_sin[10]  =  11'b11111100010;     //10pi/512
   m_cos[10]  =  11'b00111111111;     //10pi/512
   m_sin[11]  =  11'b11111011111;     //11pi/512
   m_cos[11]  =  11'b00111111110;     //11pi/512
   m_sin[12]  =  11'b11111011100;     //12pi/512
   m_cos[12]  =  11'b00111111110;     //12pi/512
   m_sin[13]  =  11'b11111011001;     //13pi/512
   m_cos[13]  =  11'b00111111110;     //13pi/512
   m_sin[14]  =  11'b11111010110;     //14pi/512
   m_cos[14]  =  11'b00111111110;     //14pi/512
   m_sin[15]  =  11'b11111010011;     //15pi/512
   m_cos[15]  =  11'b00111111110;     //15pi/512
   m_sin[16]  =  11'b11111010000;     //16pi/512
   m_cos[16]  =  11'b00111111101;     //16pi/512
   m_sin[17]  =  11'b11111001101;     //17pi/512
   m_cos[17]  =  11'b00111111101;     //17pi/512
   m_sin[18]  =  11'b11111001010;     //18pi/512
   m_cos[18]  =  11'b00111111101;     //18pi/512
   m_sin[19]  =  11'b11111000111;     //19pi/512
   m_cos[19]  =  11'b00111111100;     //19pi/512
   m_sin[20]  =  11'b11111000100;     //20pi/512
   m_cos[20]  =  11'b00111111100;     //20pi/512
   m_sin[21]  =  11'b11111000001;     //21pi/512
   m_cos[21]  =  11'b00111111100;     //21pi/512
   m_sin[22]  =  11'b11110111111;     //22pi/512
   m_cos[22]  =  11'b00111111011;     //22pi/512
   m_sin[23]  =  11'b11110111100;     //23pi/512
   m_cos[23]  =  11'b00111111011;     //23pi/512
   m_sin[24]  =  11'b11110111001;     //24pi/512
   m_cos[24]  =  11'b00111111010;     //24pi/512
   m_sin[25]  =  11'b11110110110;     //25pi/512
   m_cos[25]  =  11'b00111111010;     //25pi/512
   m_sin[26]  =  11'b11110110011;     //26pi/512
   m_cos[26]  =  11'b00111111010;     //26pi/512
   m_sin[27]  =  11'b11110110000;     //27pi/512
   m_cos[27]  =  11'b00111111001;     //27pi/512
   m_sin[28]  =  11'b11110101101;     //28pi/512
   m_cos[28]  =  11'b00111111001;     //28pi/512
   m_sin[29]  =  11'b11110101010;     //29pi/512
   m_cos[29]  =  11'b00111111000;     //29pi/512
   m_sin[30]  =  11'b11110100111;     //30pi/512
   m_cos[30]  =  11'b00111111000;     //30pi/512
   m_sin[31]  =  11'b11110100100;     //31pi/512
   m_cos[31]  =  11'b00111110111;     //31pi/512
   m_sin[32]  =  11'b11110100001;     //32pi/512
   m_cos[32]  =  11'b00111110111;     //32pi/512
   m_sin[33]  =  11'b11110011110;     //33pi/512
   m_cos[33]  =  11'b00111110110;     //33pi/512
   m_sin[34]  =  11'b11110011011;     //34pi/512
   m_cos[34]  =  11'b00111110101;     //34pi/512
   m_sin[35]  =  11'b11110011000;     //35pi/512
   m_cos[35]  =  11'b00111110101;     //35pi/512
   m_sin[36]  =  11'b11110010101;     //36pi/512
   m_cos[36]  =  11'b00111110100;     //36pi/512
   m_sin[37]  =  11'b11110010010;     //37pi/512
   m_cos[37]  =  11'b00111110100;     //37pi/512
   m_sin[38]  =  11'b11110010000;     //38pi/512
   m_cos[38]  =  11'b00111110011;     //38pi/512
   m_sin[39]  =  11'b11110001101;     //39pi/512
   m_cos[39]  =  11'b00111110010;     //39pi/512
   m_sin[40]  =  11'b11110001010;     //40pi/512
   m_cos[40]  =  11'b00111110010;     //40pi/512
   m_sin[41]  =  11'b11110000111;     //41pi/512
   m_cos[41]  =  11'b00111110001;     //41pi/512
   m_sin[42]  =  11'b11110000100;     //42pi/512
   m_cos[42]  =  11'b00111110000;     //42pi/512
   m_sin[43]  =  11'b11110000001;     //43pi/512
   m_cos[43]  =  11'b00111110000;     //43pi/512
   m_sin[44]  =  11'b11101111110;     //44pi/512
   m_cos[44]  =  11'b00111101111;     //44pi/512
   m_sin[45]  =  11'b11101111011;     //45pi/512
   m_cos[45]  =  11'b00111101110;     //45pi/512
   m_sin[46]  =  11'b11101111000;     //46pi/512
   m_cos[46]  =  11'b00111101101;     //46pi/512
   m_sin[47]  =  11'b11101110101;     //47pi/512
   m_cos[47]  =  11'b00111101100;     //47pi/512
   m_sin[48]  =  11'b11101110011;     //48pi/512
   m_cos[48]  =  11'b00111101100;     //48pi/512
   m_sin[49]  =  11'b11101110000;     //49pi/512
   m_cos[49]  =  11'b00111101011;     //49pi/512
   m_sin[50]  =  11'b11101101101;     //50pi/512
   m_cos[50]  =  11'b00111101010;     //50pi/512
   m_sin[51]  =  11'b11101101010;     //51pi/512
   m_cos[51]  =  11'b00111101001;     //51pi/512
   m_sin[52]  =  11'b11101100111;     //52pi/512
   m_cos[52]  =  11'b00111101000;     //52pi/512
   m_sin[53]  =  11'b11101100100;     //53pi/512
   m_cos[53]  =  11'b00111100111;     //53pi/512
   m_sin[54]  =  11'b11101100001;     //54pi/512
   m_cos[54]  =  11'b00111100110;     //54pi/512
   m_sin[55]  =  11'b11101011111;     //55pi/512
   m_cos[55]  =  11'b00111100101;     //55pi/512
   m_sin[56]  =  11'b11101011100;     //56pi/512
   m_cos[56]  =  11'b00111100100;     //56pi/512
   m_sin[57]  =  11'b11101011001;     //57pi/512
   m_cos[57]  =  11'b00111100011;     //57pi/512
   m_sin[58]  =  11'b11101010110;     //58pi/512
   m_cos[58]  =  11'b00111100011;     //58pi/512
   m_sin[59]  =  11'b11101010011;     //59pi/512
   m_cos[59]  =  11'b00111100010;     //59pi/512
   m_sin[60]  =  11'b11101010001;     //60pi/512
   m_cos[60]  =  11'b00111100001;     //60pi/512
   m_sin[61]  =  11'b11101001110;     //61pi/512
   m_cos[61]  =  11'b00111011111;     //61pi/512
   m_sin[62]  =  11'b11101001011;     //62pi/512
   m_cos[62]  =  11'b00111011110;     //62pi/512
   m_sin[63]  =  11'b11101001000;     //63pi/512
   m_cos[63]  =  11'b00111011101;     //63pi/512
   m_sin[64]  =  11'b11101000101;     //64pi/512
   m_cos[64]  =  11'b00111011100;     //64pi/512
   m_sin[65]  =  11'b11101000011;     //65pi/512
   m_cos[65]  =  11'b00111011011;     //65pi/512
   m_sin[66]  =  11'b11101000000;     //66pi/512
   m_cos[66]  =  11'b00111011010;     //66pi/512
   m_sin[67]  =  11'b11100111101;     //67pi/512
   m_cos[67]  =  11'b00111011001;     //67pi/512
   m_sin[68]  =  11'b11100111010;     //68pi/512
   m_cos[68]  =  11'b00111011000;     //68pi/512
   m_sin[69]  =  11'b11100111000;     //69pi/512
   m_cos[69]  =  11'b00111010111;     //69pi/512
   m_sin[70]  =  11'b11100110101;     //70pi/512
   m_cos[70]  =  11'b00111010101;     //70pi/512
   m_sin[71]  =  11'b11100110010;     //71pi/512
   m_cos[71]  =  11'b00111010100;     //71pi/512
   m_sin[72]  =  11'b11100101111;     //72pi/512
   m_cos[72]  =  11'b00111010011;     //72pi/512
   m_sin[73]  =  11'b11100101101;     //73pi/512
   m_cos[73]  =  11'b00111010010;     //73pi/512
   m_sin[74]  =  11'b11100101010;     //74pi/512
   m_cos[74]  =  11'b00111010001;     //74pi/512
   m_sin[75]  =  11'b11100100111;     //75pi/512
   m_cos[75]  =  11'b00111001111;     //75pi/512
   m_sin[76]  =  11'b11100100101;     //76pi/512
   m_cos[76]  =  11'b00111001110;     //76pi/512
   m_sin[77]  =  11'b11100100010;     //77pi/512
   m_cos[77]  =  11'b00111001101;     //77pi/512
   m_sin[78]  =  11'b11100011111;     //78pi/512
   m_cos[78]  =  11'b00111001011;     //78pi/512
   m_sin[79]  =  11'b11100011100;     //79pi/512
   m_cos[79]  =  11'b00111001010;     //79pi/512
   m_sin[80]  =  11'b11100011010;     //80pi/512
   m_cos[80]  =  11'b00111001001;     //80pi/512
   m_sin[81]  =  11'b11100010111;     //81pi/512
   m_cos[81]  =  11'b00111000111;     //81pi/512
   m_sin[82]  =  11'b11100010100;     //82pi/512
   m_cos[82]  =  11'b00111000110;     //82pi/512
   m_sin[83]  =  11'b11100010010;     //83pi/512
   m_cos[83]  =  11'b00111000101;     //83pi/512
   m_sin[84]  =  11'b11100001111;     //84pi/512
   m_cos[84]  =  11'b00111000011;     //84pi/512
   m_sin[85]  =  11'b11100001101;     //85pi/512
   m_cos[85]  =  11'b00111000010;     //85pi/512
   m_sin[86]  =  11'b11100001010;     //86pi/512
   m_cos[86]  =  11'b00111000001;     //86pi/512
   m_sin[87]  =  11'b11100000111;     //87pi/512
   m_cos[87]  =  11'b00110111111;     //87pi/512
   m_sin[88]  =  11'b11100000101;     //88pi/512
   m_cos[88]  =  11'b00110111110;     //88pi/512
   m_sin[89]  =  11'b11100000010;     //89pi/512
   m_cos[89]  =  11'b00110111100;     //89pi/512
   m_sin[90]  =  11'b11100000000;     //90pi/512
   m_cos[90]  =  11'b00110111011;     //90pi/512
   m_sin[91]  =  11'b11011111101;     //91pi/512
   m_cos[91]  =  11'b00110111001;     //91pi/512
   m_sin[92]  =  11'b11011111010;     //92pi/512
   m_cos[92]  =  11'b00110111000;     //92pi/512
   m_sin[93]  =  11'b11011111000;     //93pi/512
   m_cos[93]  =  11'b00110110110;     //93pi/512
   m_sin[94]  =  11'b11011110101;     //94pi/512
   m_cos[94]  =  11'b00110110101;     //94pi/512
   m_sin[95]  =  11'b11011110011;     //95pi/512
   m_cos[95]  =  11'b00110110011;     //95pi/512
   m_sin[96]  =  11'b11011110000;     //96pi/512
   m_cos[96]  =  11'b00110110001;     //96pi/512
   m_sin[97]  =  11'b11011101110;     //97pi/512
   m_cos[97]  =  11'b00110110000;     //97pi/512
   m_sin[98]  =  11'b11011101011;     //98pi/512
   m_cos[98]  =  11'b00110101110;     //98pi/512
   m_sin[99]  =  11'b11011101001;     //99pi/512
   m_cos[99]  =  11'b00110101101;     //99pi/512
   m_sin[100]  =  11'b11011100110;     //100pi/512
   m_cos[100]  =  11'b00110101011;     //100pi/512
   m_sin[101]  =  11'b11011100100;     //101pi/512
   m_cos[101]  =  11'b00110101001;     //101pi/512
   m_sin[102]  =  11'b11011100001;     //102pi/512
   m_cos[102]  =  11'b00110101000;     //102pi/512
   m_sin[103]  =  11'b11011011111;     //103pi/512
   m_cos[103]  =  11'b00110100110;     //103pi/512
   m_sin[104]  =  11'b11011011100;     //104pi/512
   m_cos[104]  =  11'b00110100100;     //104pi/512
   m_sin[105]  =  11'b11011011010;     //105pi/512
   m_cos[105]  =  11'b00110100011;     //105pi/512
   m_sin[106]  =  11'b11011010111;     //106pi/512
   m_cos[106]  =  11'b00110100001;     //106pi/512
   m_sin[107]  =  11'b11011010101;     //107pi/512
   m_cos[107]  =  11'b00110011111;     //107pi/512
   m_sin[108]  =  11'b11011010011;     //108pi/512
   m_cos[108]  =  11'b00110011101;     //108pi/512
   m_sin[109]  =  11'b11011010000;     //109pi/512
   m_cos[109]  =  11'b00110011100;     //109pi/512
   m_sin[110]  =  11'b11011001110;     //110pi/512
   m_cos[110]  =  11'b00110011010;     //110pi/512
   m_sin[111]  =  11'b11011001011;     //111pi/512
   m_cos[111]  =  11'b00110011000;     //111pi/512
   m_sin[112]  =  11'b11011001001;     //112pi/512
   m_cos[112]  =  11'b00110010110;     //112pi/512
   m_sin[113]  =  11'b11011000111;     //113pi/512
   m_cos[113]  =  11'b00110010100;     //113pi/512
   m_sin[114]  =  11'b11011000100;     //114pi/512
   m_cos[114]  =  11'b00110010011;     //114pi/512
   m_sin[115]  =  11'b11011000010;     //115pi/512
   m_cos[115]  =  11'b00110010001;     //115pi/512
   m_sin[116]  =  11'b11011000000;     //116pi/512
   m_cos[116]  =  11'b00110001111;     //116pi/512
   m_sin[117]  =  11'b11010111101;     //117pi/512
   m_cos[117]  =  11'b00110001101;     //117pi/512
   m_sin[118]  =  11'b11010111011;     //118pi/512
   m_cos[118]  =  11'b00110001011;     //118pi/512
   m_sin[119]  =  11'b11010111001;     //119pi/512
   m_cos[119]  =  11'b00110001001;     //119pi/512
   m_sin[120]  =  11'b11010110110;     //120pi/512
   m_cos[120]  =  11'b00110000111;     //120pi/512
   m_sin[121]  =  11'b11010110100;     //121pi/512
   m_cos[121]  =  11'b00110000101;     //121pi/512
   m_sin[122]  =  11'b11010110010;     //122pi/512
   m_cos[122]  =  11'b00110000011;     //122pi/512
   m_sin[123]  =  11'b11010110000;     //123pi/512
   m_cos[123]  =  11'b00110000001;     //123pi/512
   m_sin[124]  =  11'b11010101101;     //124pi/512
   m_cos[124]  =  11'b00101111111;     //124pi/512
   m_sin[125]  =  11'b11010101011;     //125pi/512
   m_cos[125]  =  11'b00101111101;     //125pi/512
   m_sin[126]  =  11'b11010101001;     //126pi/512
   m_cos[126]  =  11'b00101111011;     //126pi/512
   m_sin[127]  =  11'b11010100111;     //127pi/512
   m_cos[127]  =  11'b00101111001;     //127pi/512
   m_sin[128]  =  11'b11010100100;     //128pi/512
   m_cos[128]  =  11'b00101110111;     //128pi/512
   m_sin[129]  =  11'b11010100010;     //129pi/512
   m_cos[129]  =  11'b00101110101;     //129pi/512
   m_sin[130]  =  11'b11010100000;     //130pi/512
   m_cos[130]  =  11'b00101110011;     //130pi/512
   m_sin[131]  =  11'b11010011110;     //131pi/512
   m_cos[131]  =  11'b00101110001;     //131pi/512
   m_sin[132]  =  11'b11010011100;     //132pi/512
   m_cos[132]  =  11'b00101101111;     //132pi/512
   m_sin[133]  =  11'b11010011010;     //133pi/512
   m_cos[133]  =  11'b00101101101;     //133pi/512
   m_sin[134]  =  11'b11010011000;     //134pi/512
   m_cos[134]  =  11'b00101101011;     //134pi/512
   m_sin[135]  =  11'b11010010101;     //135pi/512
   m_cos[135]  =  11'b00101101001;     //135pi/512
   m_sin[136]  =  11'b11010010011;     //136pi/512
   m_cos[136]  =  11'b00101100111;     //136pi/512
   m_sin[137]  =  11'b11010010001;     //137pi/512
   m_cos[137]  =  11'b00101100101;     //137pi/512
   m_sin[138]  =  11'b11010001111;     //138pi/512
   m_cos[138]  =  11'b00101100011;     //138pi/512
   m_sin[139]  =  11'b11010001101;     //139pi/512
   m_cos[139]  =  11'b00101100000;     //139pi/512
   m_sin[140]  =  11'b11010001011;     //140pi/512
   m_cos[140]  =  11'b00101011110;     //140pi/512
   m_sin[141]  =  11'b11010001001;     //141pi/512
   m_cos[141]  =  11'b00101011100;     //141pi/512
   m_sin[142]  =  11'b11010000111;     //142pi/512
   m_cos[142]  =  11'b00101011010;     //142pi/512
   m_sin[143]  =  11'b11010000101;     //143pi/512
   m_cos[143]  =  11'b00101011000;     //143pi/512
   m_sin[144]  =  11'b11010000011;     //144pi/512
   m_cos[144]  =  11'b00101010101;     //144pi/512
   m_sin[145]  =  11'b11010000001;     //145pi/512
   m_cos[145]  =  11'b00101010011;     //145pi/512
   m_sin[146]  =  11'b11001111111;     //146pi/512
   m_cos[146]  =  11'b00101010001;     //146pi/512
   m_sin[147]  =  11'b11001111101;     //147pi/512
   m_cos[147]  =  11'b00101001111;     //147pi/512
   m_sin[148]  =  11'b11001111011;     //148pi/512
   m_cos[148]  =  11'b00101001100;     //148pi/512
   m_sin[149]  =  11'b11001111001;     //149pi/512
   m_cos[149]  =  11'b00101001010;     //149pi/512
   m_sin[150]  =  11'b11001110111;     //150pi/512
   m_cos[150]  =  11'b00101001000;     //150pi/512
   m_sin[151]  =  11'b11001110101;     //151pi/512
   m_cos[151]  =  11'b00101000110;     //151pi/512
   m_sin[152]  =  11'b11001110011;     //152pi/512
   m_cos[152]  =  11'b00101000011;     //152pi/512
   m_sin[153]  =  11'b11001110010;     //153pi/512
   m_cos[153]  =  11'b00101000001;     //153pi/512
   m_sin[154]  =  11'b11001110000;     //154pi/512
   m_cos[154]  =  11'b00100111111;     //154pi/512
   m_sin[155]  =  11'b11001101110;     //155pi/512
   m_cos[155]  =  11'b00100111100;     //155pi/512
   m_sin[156]  =  11'b11001101100;     //156pi/512
   m_cos[156]  =  11'b00100111010;     //156pi/512
   m_sin[157]  =  11'b11001101010;     //157pi/512
   m_cos[157]  =  11'b00100111000;     //157pi/512
   m_sin[158]  =  11'b11001101000;     //158pi/512
   m_cos[158]  =  11'b00100110101;     //158pi/512
   m_sin[159]  =  11'b11001100111;     //159pi/512
   m_cos[159]  =  11'b00100110011;     //159pi/512
   m_sin[160]  =  11'b11001100101;     //160pi/512
   m_cos[160]  =  11'b00100110000;     //160pi/512
   m_sin[161]  =  11'b11001100011;     //161pi/512
   m_cos[161]  =  11'b00100101110;     //161pi/512
   m_sin[162]  =  11'b11001100001;     //162pi/512
   m_cos[162]  =  11'b00100101100;     //162pi/512
   m_sin[163]  =  11'b11001011111;     //163pi/512
   m_cos[163]  =  11'b00100101001;     //163pi/512
   m_sin[164]  =  11'b11001011110;     //164pi/512
   m_cos[164]  =  11'b00100100111;     //164pi/512
   m_sin[165]  =  11'b11001011100;     //165pi/512
   m_cos[165]  =  11'b00100100100;     //165pi/512
   m_sin[166]  =  11'b11001011010;     //166pi/512
   m_cos[166]  =  11'b00100100010;     //166pi/512
   m_sin[167]  =  11'b11001011001;     //167pi/512
   m_cos[167]  =  11'b00100011111;     //167pi/512
   m_sin[168]  =  11'b11001010111;     //168pi/512
   m_cos[168]  =  11'b00100011101;     //168pi/512
   m_sin[169]  =  11'b11001010101;     //169pi/512
   m_cos[169]  =  11'b00100011011;     //169pi/512
   m_sin[170]  =  11'b11001010100;     //170pi/512
   m_cos[170]  =  11'b00100011000;     //170pi/512
   m_sin[171]  =  11'b11001010010;     //171pi/512
   m_cos[171]  =  11'b00100010110;     //171pi/512
   m_sin[172]  =  11'b11001010000;     //172pi/512
   m_cos[172]  =  11'b00100010011;     //172pi/512
   m_sin[173]  =  11'b11001001111;     //173pi/512
   m_cos[173]  =  11'b00100010000;     //173pi/512
   m_sin[174]  =  11'b11001001101;     //174pi/512
   m_cos[174]  =  11'b00100001110;     //174pi/512
   m_sin[175]  =  11'b11001001100;     //175pi/512
   m_cos[175]  =  11'b00100001011;     //175pi/512
   m_sin[176]  =  11'b11001001010;     //176pi/512
   m_cos[176]  =  11'b00100001001;     //176pi/512
   m_sin[177]  =  11'b11001001001;     //177pi/512
   m_cos[177]  =  11'b00100000110;     //177pi/512
   m_sin[178]  =  11'b11001000111;     //178pi/512
   m_cos[178]  =  11'b00100000100;     //178pi/512
   m_sin[179]  =  11'b11001000110;     //179pi/512
   m_cos[179]  =  11'b00100000001;     //179pi/512
   m_sin[180]  =  11'b11001000100;     //180pi/512
   m_cos[180]  =  11'b00011111111;     //180pi/512
   m_sin[181]  =  11'b11001000011;     //181pi/512
   m_cos[181]  =  11'b00011111100;     //181pi/512
   m_sin[182]  =  11'b11001000001;     //182pi/512
   m_cos[182]  =  11'b00011111001;     //182pi/512
   m_sin[183]  =  11'b11001000000;     //183pi/512
   m_cos[183]  =  11'b00011110111;     //183pi/512
   m_sin[184]  =  11'b11000111110;     //184pi/512
   m_cos[184]  =  11'b00011110100;     //184pi/512
   m_sin[185]  =  11'b11000111101;     //185pi/512
   m_cos[185]  =  11'b00011110010;     //185pi/512
   m_sin[186]  =  11'b11000111011;     //186pi/512
   m_cos[186]  =  11'b00011101111;     //186pi/512
   m_sin[187]  =  11'b11000111010;     //187pi/512
   m_cos[187]  =  11'b00011101100;     //187pi/512
   m_sin[188]  =  11'b11000111001;     //188pi/512
   m_cos[188]  =  11'b00011101010;     //188pi/512
   m_sin[189]  =  11'b11000110111;     //189pi/512
   m_cos[189]  =  11'b00011100111;     //189pi/512
   m_sin[190]  =  11'b11000110110;     //190pi/512
   m_cos[190]  =  11'b00011100100;     //190pi/512
   m_sin[191]  =  11'b11000110101;     //191pi/512
   m_cos[191]  =  11'b00011100010;     //191pi/512
   m_sin[192]  =  11'b11000110011;     //192pi/512
   m_cos[192]  =  11'b00011011111;     //192pi/512
   m_sin[193]  =  11'b11000110010;     //193pi/512
   m_cos[193]  =  11'b00011011100;     //193pi/512
   m_sin[194]  =  11'b11000110001;     //194pi/512
   m_cos[194]  =  11'b00011011010;     //194pi/512
   m_sin[195]  =  11'b11000101111;     //195pi/512
   m_cos[195]  =  11'b00011010111;     //195pi/512
   m_sin[196]  =  11'b11000101110;     //196pi/512
   m_cos[196]  =  11'b00011010100;     //196pi/512
   m_sin[197]  =  11'b11000101101;     //197pi/512
   m_cos[197]  =  11'b00011010001;     //197pi/512
   m_sin[198]  =  11'b11000101100;     //198pi/512
   m_cos[198]  =  11'b00011001111;     //198pi/512
   m_sin[199]  =  11'b11000101011;     //199pi/512
   m_cos[199]  =  11'b00011001100;     //199pi/512
   m_sin[200]  =  11'b11000101001;     //200pi/512
   m_cos[200]  =  11'b00011001001;     //200pi/512
   m_sin[201]  =  11'b11000101000;     //201pi/512
   m_cos[201]  =  11'b00011000110;     //201pi/512
   m_sin[202]  =  11'b11000100111;     //202pi/512
   m_cos[202]  =  11'b00011000100;     //202pi/512
   m_sin[203]  =  11'b11000100110;     //203pi/512
   m_cos[203]  =  11'b00011000001;     //203pi/512
   m_sin[204]  =  11'b11000100101;     //204pi/512
   m_cos[204]  =  11'b00010111110;     //204pi/512
   m_sin[205]  =  11'b11000100100;     //205pi/512
   m_cos[205]  =  11'b00010111011;     //205pi/512
   m_sin[206]  =  11'b11000100011;     //206pi/512
   m_cos[206]  =  11'b00010111001;     //206pi/512
   m_sin[207]  =  11'b11000100010;     //207pi/512
   m_cos[207]  =  11'b00010110110;     //207pi/512
   m_sin[208]  =  11'b11000100001;     //208pi/512
   m_cos[208]  =  11'b00010110011;     //208pi/512
   m_sin[209]  =  11'b11000011111;     //209pi/512
   m_cos[209]  =  11'b00010110000;     //209pi/512
   m_sin[210]  =  11'b11000011110;     //210pi/512
   m_cos[210]  =  11'b00010101101;     //210pi/512
   m_sin[211]  =  11'b11000011101;     //211pi/512
   m_cos[211]  =  11'b00010101011;     //211pi/512
   m_sin[212]  =  11'b11000011100;     //212pi/512
   m_cos[212]  =  11'b00010101000;     //212pi/512
   m_sin[213]  =  11'b11000011011;     //213pi/512
   m_cos[213]  =  11'b00010100101;     //213pi/512
   m_sin[214]  =  11'b11000011011;     //214pi/512
   m_cos[214]  =  11'b00010100010;     //214pi/512
   m_sin[215]  =  11'b11000011010;     //215pi/512
   m_cos[215]  =  11'b00010011111;     //215pi/512
   m_sin[216]  =  11'b11000011001;     //216pi/512
   m_cos[216]  =  11'b00010011101;     //216pi/512
   m_sin[217]  =  11'b11000011000;     //217pi/512
   m_cos[217]  =  11'b00010011010;     //217pi/512
   m_sin[218]  =  11'b11000010111;     //218pi/512
   m_cos[218]  =  11'b00010010111;     //218pi/512
   m_sin[219]  =  11'b11000010110;     //219pi/512
   m_cos[219]  =  11'b00010010100;     //219pi/512
   m_sin[220]  =  11'b11000010101;     //220pi/512
   m_cos[220]  =  11'b00010010001;     //220pi/512
   m_sin[221]  =  11'b11000010100;     //221pi/512
   m_cos[221]  =  11'b00010001110;     //221pi/512
   m_sin[222]  =  11'b11000010011;     //222pi/512
   m_cos[222]  =  11'b00010001011;     //222pi/512
   m_sin[223]  =  11'b11000010011;     //223pi/512
   m_cos[223]  =  11'b00010001001;     //223pi/512
   m_sin[224]  =  11'b11000010010;     //224pi/512
   m_cos[224]  =  11'b00010000110;     //224pi/512
   m_sin[225]  =  11'b11000010001;     //225pi/512
   m_cos[225]  =  11'b00010000011;     //225pi/512
   m_sin[226]  =  11'b11000010000;     //226pi/512
   m_cos[226]  =  11'b00010000000;     //226pi/512
   m_sin[227]  =  11'b11000010000;     //227pi/512
   m_cos[227]  =  11'b00001111101;     //227pi/512
   m_sin[228]  =  11'b11000001111;     //228pi/512
   m_cos[228]  =  11'b00001111010;     //228pi/512
   m_sin[229]  =  11'b11000001110;     //229pi/512
   m_cos[229]  =  11'b00001110111;     //229pi/512
   m_sin[230]  =  11'b11000001101;     //230pi/512
   m_cos[230]  =  11'b00001110100;     //230pi/512
   m_sin[231]  =  11'b11000001101;     //231pi/512
   m_cos[231]  =  11'b00001110001;     //231pi/512
   m_sin[232]  =  11'b11000001100;     //232pi/512
   m_cos[232]  =  11'b00001101110;     //232pi/512
   m_sin[233]  =  11'b11000001100;     //233pi/512
   m_cos[233]  =  11'b00001101100;     //233pi/512
   m_sin[234]  =  11'b11000001011;     //234pi/512
   m_cos[234]  =  11'b00001101001;     //234pi/512
   m_sin[235]  =  11'b11000001010;     //235pi/512
   m_cos[235]  =  11'b00001100110;     //235pi/512
   m_sin[236]  =  11'b11000001010;     //236pi/512
   m_cos[236]  =  11'b00001100011;     //236pi/512
   m_sin[237]  =  11'b11000001001;     //237pi/512
   m_cos[237]  =  11'b00001100000;     //237pi/512
   m_sin[238]  =  11'b11000001001;     //238pi/512
   m_cos[238]  =  11'b00001011101;     //238pi/512
   m_sin[239]  =  11'b11000001000;     //239pi/512
   m_cos[239]  =  11'b00001011010;     //239pi/512
   m_sin[240]  =  11'b11000001000;     //240pi/512
   m_cos[240]  =  11'b00001010111;     //240pi/512
   m_sin[241]  =  11'b11000000111;     //241pi/512
   m_cos[241]  =  11'b00001010100;     //241pi/512
   m_sin[242]  =  11'b11000000111;     //242pi/512
   m_cos[242]  =  11'b00001010001;     //242pi/512
   m_sin[243]  =  11'b11000000110;     //243pi/512
   m_cos[243]  =  11'b00001001110;     //243pi/512
   m_sin[244]  =  11'b11000000110;     //244pi/512
   m_cos[244]  =  11'b00001001011;     //244pi/512
   m_sin[245]  =  11'b11000000101;     //245pi/512
   m_cos[245]  =  11'b00001001000;     //245pi/512
   m_sin[246]  =  11'b11000000101;     //246pi/512
   m_cos[246]  =  11'b00001000101;     //246pi/512
   m_sin[247]  =  11'b11000000100;     //247pi/512
   m_cos[247]  =  11'b00001000010;     //247pi/512
   m_sin[248]  =  11'b11000000100;     //248pi/512
   m_cos[248]  =  11'b00000111111;     //248pi/512
   m_sin[249]  =  11'b11000000100;     //249pi/512
   m_cos[249]  =  11'b00000111100;     //249pi/512
   m_sin[250]  =  11'b11000000011;     //250pi/512
   m_cos[250]  =  11'b00000111001;     //250pi/512
   m_sin[251]  =  11'b11000000011;     //251pi/512
   m_cos[251]  =  11'b00000110111;     //251pi/512
   m_sin[252]  =  11'b11000000011;     //252pi/512
   m_cos[252]  =  11'b00000110100;     //252pi/512
   m_sin[253]  =  11'b11000000010;     //253pi/512
   m_cos[253]  =  11'b00000110001;     //253pi/512
   m_sin[254]  =  11'b11000000010;     //254pi/512
   m_cos[254]  =  11'b00000101110;     //254pi/512
   m_sin[255]  =  11'b11000000010;     //255pi/512
   m_cos[255]  =  11'b00000101011;     //255pi/512
   m_sin[256]  =  11'b11000000010;     //256pi/512
   m_cos[256]  =  11'b00000101000;     //256pi/512
   m_sin[257]  =  11'b11000000001;     //257pi/512
   m_cos[257]  =  11'b00000100101;     //257pi/512
   m_sin[258]  =  11'b11000000001;     //258pi/512
   m_cos[258]  =  11'b00000100010;     //258pi/512
   m_sin[259]  =  11'b11000000001;     //259pi/512
   m_cos[259]  =  11'b00000011111;     //259pi/512
   m_sin[260]  =  11'b11000000001;     //260pi/512
   m_cos[260]  =  11'b00000011100;     //260pi/512
   m_sin[261]  =  11'b11000000001;     //261pi/512
   m_cos[261]  =  11'b00000011001;     //261pi/512
   m_sin[262]  =  11'b11000000000;     //262pi/512
   m_cos[262]  =  11'b00000010110;     //262pi/512
   m_sin[263]  =  11'b11000000000;     //263pi/512
   m_cos[263]  =  11'b00000010011;     //263pi/512
   m_sin[264]  =  11'b11000000000;     //264pi/512
   m_cos[264]  =  11'b00000010000;     //264pi/512
   m_sin[265]  =  11'b11000000000;     //265pi/512
   m_cos[265]  =  11'b00000001101;     //265pi/512
   m_sin[266]  =  11'b11000000000;     //266pi/512
   m_cos[266]  =  11'b00000001010;     //266pi/512
   m_sin[267]  =  11'b11000000000;     //267pi/512
   m_cos[267]  =  11'b00000000111;     //267pi/512
   m_sin[268]  =  11'b11000000000;     //268pi/512
   m_cos[268]  =  11'b00000000100;     //268pi/512
   m_sin[269]  =  11'b11000000000;     //269pi/512
   m_cos[269]  =  11'b00000000001;     //269pi/512
   m_sin[270]  =  11'b11000000000;     //270pi/512
   m_cos[270]  =  11'b11111111110;     //270pi/512
   m_sin[271]  =  11'b11000000000;     //271pi/512
   m_cos[271]  =  11'b11111111011;     //271pi/512
   m_sin[272]  =  11'b11000000000;     //272pi/512
   m_cos[272]  =  11'b11111111000;     //272pi/512
   m_sin[273]  =  11'b11000000000;     //273pi/512
   m_cos[273]  =  11'b11111110101;     //273pi/512
   m_sin[274]  =  11'b11000000000;     //274pi/512
   m_cos[274]  =  11'b11111110010;     //274pi/512
   m_sin[275]  =  11'b11000000000;     //275pi/512
   m_cos[275]  =  11'b11111110000;     //275pi/512
   m_sin[276]  =  11'b11000000000;     //276pi/512
   m_cos[276]  =  11'b11111101101;     //276pi/512
   m_sin[277]  =  11'b11000000000;     //277pi/512
   m_cos[277]  =  11'b11111101010;     //277pi/512
   m_sin[278]  =  11'b11000000001;     //278pi/512
   m_cos[278]  =  11'b11111100111;     //278pi/512
   m_sin[279]  =  11'b11000000001;     //279pi/512
   m_cos[279]  =  11'b11111100100;     //279pi/512
   m_sin[280]  =  11'b11000000001;     //280pi/512
   m_cos[280]  =  11'b11111100001;     //280pi/512
   m_sin[281]  =  11'b11000000001;     //281pi/512
   m_cos[281]  =  11'b11111011110;     //281pi/512
   m_sin[282]  =  11'b11000000001;     //282pi/512
   m_cos[282]  =  11'b11111011011;     //282pi/512
   m_sin[283]  =  11'b11000000010;     //283pi/512
   m_cos[283]  =  11'b11111011000;     //283pi/512
   m_sin[284]  =  11'b11000000010;     //284pi/512
   m_cos[284]  =  11'b11111010101;     //284pi/512
   m_sin[285]  =  11'b11000000010;     //285pi/512
   m_cos[285]  =  11'b11111010010;     //285pi/512
   m_sin[286]  =  11'b11000000010;     //286pi/512
   m_cos[286]  =  11'b11111001111;     //286pi/512
   m_sin[287]  =  11'b11000000011;     //287pi/512
   m_cos[287]  =  11'b11111001100;     //287pi/512
   m_sin[288]  =  11'b11000000011;     //288pi/512
   m_cos[288]  =  11'b11111001001;     //288pi/512
   m_sin[289]  =  11'b11000000011;     //289pi/512
   m_cos[289]  =  11'b11111000110;     //289pi/512
   m_sin[290]  =  11'b11000000100;     //290pi/512
   m_cos[290]  =  11'b11111000011;     //290pi/512
   m_sin[291]  =  11'b11000000100;     //291pi/512
   m_cos[291]  =  11'b11111000000;     //291pi/512
   m_sin[292]  =  11'b11000000100;     //292pi/512
   m_cos[292]  =  11'b11110111101;     //292pi/512
   m_sin[293]  =  11'b11000000101;     //293pi/512
   m_cos[293]  =  11'b11110111010;     //293pi/512
   m_sin[294]  =  11'b11000000101;     //294pi/512
   m_cos[294]  =  11'b11110110111;     //294pi/512
   m_sin[295]  =  11'b11000000110;     //295pi/512
   m_cos[295]  =  11'b11110110100;     //295pi/512
   m_sin[296]  =  11'b11000000110;     //296pi/512
   m_cos[296]  =  11'b11110110001;     //296pi/512
   m_sin[297]  =  11'b11000000111;     //297pi/512
   m_cos[297]  =  11'b11110101110;     //297pi/512
   m_sin[298]  =  11'b11000000111;     //298pi/512
   m_cos[298]  =  11'b11110101011;     //298pi/512
   m_sin[299]  =  11'b11000001000;     //299pi/512
   m_cos[299]  =  11'b11110101000;     //299pi/512
   m_sin[300]  =  11'b11000001000;     //300pi/512
   m_cos[300]  =  11'b11110100101;     //300pi/512
   m_sin[301]  =  11'b11000001001;     //301pi/512
   m_cos[301]  =  11'b11110100010;     //301pi/512
   m_sin[302]  =  11'b11000001001;     //302pi/512
   m_cos[302]  =  11'b11110100000;     //302pi/512
   m_sin[303]  =  11'b11000001010;     //303pi/512
   m_cos[303]  =  11'b11110011101;     //303pi/512
   m_sin[304]  =  11'b11000001010;     //304pi/512
   m_cos[304]  =  11'b11110011010;     //304pi/512
   m_sin[305]  =  11'b11000001011;     //305pi/512
   m_cos[305]  =  11'b11110010111;     //305pi/512
   m_sin[306]  =  11'b11000001100;     //306pi/512
   m_cos[306]  =  11'b11110010100;     //306pi/512
   m_sin[307]  =  11'b11000001100;     //307pi/512
   m_cos[307]  =  11'b11110010001;     //307pi/512
   m_sin[308]  =  11'b11000001101;     //308pi/512
   m_cos[308]  =  11'b11110001110;     //308pi/512
   m_sin[309]  =  11'b11000001110;     //309pi/512
   m_cos[309]  =  11'b11110001011;     //309pi/512
   m_sin[310]  =  11'b11000001110;     //310pi/512
   m_cos[310]  =  11'b11110001000;     //310pi/512
   m_sin[311]  =  11'b11000001111;     //311pi/512
   m_cos[311]  =  11'b11110000101;     //311pi/512
   m_sin[312]  =  11'b11000010000;     //312pi/512
   m_cos[312]  =  11'b11110000010;     //312pi/512
   m_sin[313]  =  11'b11000010000;     //313pi/512
   m_cos[313]  =  11'b11101111111;     //313pi/512
   m_sin[314]  =  11'b11000010001;     //314pi/512
   m_cos[314]  =  11'b11101111101;     //314pi/512
   m_sin[315]  =  11'b11000010010;     //315pi/512
   m_cos[315]  =  11'b11101111010;     //315pi/512
   m_sin[316]  =  11'b11000010011;     //316pi/512
   m_cos[316]  =  11'b11101110111;     //316pi/512
   m_sin[317]  =  11'b11000010100;     //317pi/512
   m_cos[317]  =  11'b11101110100;     //317pi/512
   m_sin[318]  =  11'b11000010100;     //318pi/512
   m_cos[318]  =  11'b11101110001;     //318pi/512
   m_sin[319]  =  11'b11000010101;     //319pi/512
   m_cos[319]  =  11'b11101101110;     //319pi/512
   m_sin[320]  =  11'b11000010110;     //320pi/512
   m_cos[320]  =  11'b11101101011;     //320pi/512
   m_sin[321]  =  11'b11000010111;     //321pi/512
   m_cos[321]  =  11'b11101101001;     //321pi/512
   m_sin[322]  =  11'b11000011000;     //322pi/512
   m_cos[322]  =  11'b11101100110;     //322pi/512
   m_sin[323]  =  11'b11000011001;     //323pi/512
   m_cos[323]  =  11'b11101100011;     //323pi/512
   m_sin[324]  =  11'b11000011010;     //324pi/512
   m_cos[324]  =  11'b11101100000;     //324pi/512
   m_sin[325]  =  11'b11000011011;     //325pi/512
   m_cos[325]  =  11'b11101011101;     //325pi/512
   m_sin[326]  =  11'b11000011100;     //326pi/512
   m_cos[326]  =  11'b11101011010;     //326pi/512
   m_sin[327]  =  11'b11000011101;     //327pi/512
   m_cos[327]  =  11'b11101011000;     //327pi/512
   m_sin[328]  =  11'b11000011110;     //328pi/512
   m_cos[328]  =  11'b11101010101;     //328pi/512
   m_sin[329]  =  11'b11000011111;     //329pi/512
   m_cos[329]  =  11'b11101010010;     //329pi/512
   m_sin[330]  =  11'b11000100000;     //330pi/512
   m_cos[330]  =  11'b11101001111;     //330pi/512
   m_sin[331]  =  11'b11000100001;     //331pi/512
   m_cos[331]  =  11'b11101001100;     //331pi/512
   m_sin[332]  =  11'b11000100010;     //332pi/512
   m_cos[332]  =  11'b11101001001;     //332pi/512
   m_sin[333]  =  11'b11000100011;     //333pi/512
   m_cos[333]  =  11'b11101000111;     //333pi/512
   m_sin[334]  =  11'b11000100100;     //334pi/512
   m_cos[334]  =  11'b11101000100;     //334pi/512
   m_sin[335]  =  11'b11000100101;     //335pi/512
   m_cos[335]  =  11'b11101000001;     //335pi/512
   m_sin[336]  =  11'b11000100110;     //336pi/512
   m_cos[336]  =  11'b11100111110;     //336pi/512
   m_sin[337]  =  11'b11000100111;     //337pi/512
   m_cos[337]  =  11'b11100111100;     //337pi/512
   m_sin[338]  =  11'b11000101000;     //338pi/512
   m_cos[338]  =  11'b11100111001;     //338pi/512
   m_sin[339]  =  11'b11000101001;     //339pi/512
   m_cos[339]  =  11'b11100110110;     //339pi/512
   m_sin[340]  =  11'b11000101011;     //340pi/512
   m_cos[340]  =  11'b11100110011;     //340pi/512
   m_sin[341]  =  11'b11000101100;     //341pi/512
   m_cos[341]  =  11'b11100110001;     //341pi/512
   m_sin[342]  =  11'b11000101101;     //342pi/512
   m_cos[342]  =  11'b11100101110;     //342pi/512
   m_sin[343]  =  11'b11000101110;     //343pi/512
   m_cos[343]  =  11'b11100101011;     //343pi/512
   m_sin[344]  =  11'b11000110000;     //344pi/512
   m_cos[344]  =  11'b11100101001;     //344pi/512
   m_sin[345]  =  11'b11000110001;     //345pi/512
   m_cos[345]  =  11'b11100100110;     //345pi/512
   m_sin[346]  =  11'b11000110010;     //346pi/512
   m_cos[346]  =  11'b11100100011;     //346pi/512
   m_sin[347]  =  11'b11000110011;     //347pi/512
   m_cos[347]  =  11'b11100100000;     //347pi/512
   m_sin[348]  =  11'b11000110101;     //348pi/512
   m_cos[348]  =  11'b11100011110;     //348pi/512
   m_sin[349]  =  11'b11000110110;     //349pi/512
   m_cos[349]  =  11'b11100011011;     //349pi/512
   m_sin[350]  =  11'b11000110111;     //350pi/512
   m_cos[350]  =  11'b11100011000;     //350pi/512
   m_sin[351]  =  11'b11000111001;     //351pi/512
   m_cos[351]  =  11'b11100010110;     //351pi/512
   m_sin[352]  =  11'b11000111010;     //352pi/512
   m_cos[352]  =  11'b11100010011;     //352pi/512
   m_sin[353]  =  11'b11000111011;     //353pi/512
   m_cos[353]  =  11'b11100010000;     //353pi/512
   m_sin[354]  =  11'b11000111101;     //354pi/512
   m_cos[354]  =  11'b11100001110;     //354pi/512
   m_sin[355]  =  11'b11000111110;     //355pi/512
   m_cos[355]  =  11'b11100001011;     //355pi/512
   m_sin[356]  =  11'b11001000000;     //356pi/512
   m_cos[356]  =  11'b11100001001;     //356pi/512
   m_sin[357]  =  11'b11001000001;     //357pi/512
   m_cos[357]  =  11'b11100000110;     //357pi/512
   m_sin[358]  =  11'b11001000011;     //358pi/512
   m_cos[358]  =  11'b11100000011;     //358pi/512
   m_sin[359]  =  11'b11001000100;     //359pi/512
   m_cos[359]  =  11'b11100000001;     //359pi/512
   m_sin[360]  =  11'b11001000110;     //360pi/512
   m_cos[360]  =  11'b11011111110;     //360pi/512
   m_sin[361]  =  11'b11001000111;     //361pi/512
   m_cos[361]  =  11'b11011111100;     //361pi/512
   m_sin[362]  =  11'b11001001001;     //362pi/512
   m_cos[362]  =  11'b11011111001;     //362pi/512
   m_sin[363]  =  11'b11001001010;     //363pi/512
   m_cos[363]  =  11'b11011110110;     //363pi/512
   m_sin[364]  =  11'b11001001100;     //364pi/512
   m_cos[364]  =  11'b11011110100;     //364pi/512
   m_sin[365]  =  11'b11001001101;     //365pi/512
   m_cos[365]  =  11'b11011110001;     //365pi/512
   m_sin[366]  =  11'b11001001111;     //366pi/512
   m_cos[366]  =  11'b11011101111;     //366pi/512
   m_sin[367]  =  11'b11001010001;     //367pi/512
   m_cos[367]  =  11'b11011101100;     //367pi/512
   m_sin[368]  =  11'b11001010010;     //368pi/512
   m_cos[368]  =  11'b11011101010;     //368pi/512
   m_sin[369]  =  11'b11001010100;     //369pi/512
   m_cos[369]  =  11'b11011100111;     //369pi/512
   m_sin[370]  =  11'b11001010101;     //370pi/512
   m_cos[370]  =  11'b11011100101;     //370pi/512
   m_sin[371]  =  11'b11001010111;     //371pi/512
   m_cos[371]  =  11'b11011100010;     //371pi/512
   m_sin[372]  =  11'b11001011001;     //372pi/512
   m_cos[372]  =  11'b11011100000;     //372pi/512
   m_sin[373]  =  11'b11001011010;     //373pi/512
   m_cos[373]  =  11'b11011011101;     //373pi/512
   m_sin[374]  =  11'b11001011100;     //374pi/512
   m_cos[374]  =  11'b11011011011;     //374pi/512
   m_sin[375]  =  11'b11001011110;     //375pi/512
   m_cos[375]  =  11'b11011011001;     //375pi/512
   m_sin[376]  =  11'b11001100000;     //376pi/512
   m_cos[376]  =  11'b11011010110;     //376pi/512
   m_sin[377]  =  11'b11001100001;     //377pi/512
   m_cos[377]  =  11'b11011010100;     //377pi/512
   m_sin[378]  =  11'b11001100011;     //378pi/512
   m_cos[378]  =  11'b11011010001;     //378pi/512
   m_sin[379]  =  11'b11001100101;     //379pi/512
   m_cos[379]  =  11'b11011001111;     //379pi/512
   m_sin[380]  =  11'b11001100111;     //380pi/512
   m_cos[380]  =  11'b11011001100;     //380pi/512
   m_sin[381]  =  11'b11001101000;     //381pi/512
   m_cos[381]  =  11'b11011001010;     //381pi/512
   m_sin[382]  =  11'b11001101010;     //382pi/512
   m_cos[382]  =  11'b11011001000;     //382pi/512
   m_sin[383]  =  11'b11001101100;     //383pi/512
   m_cos[383]  =  11'b11011000101;     //383pi/512
   m_sin[384]  =  11'b11001101110;     //384pi/512
   m_cos[384]  =  11'b11011000011;     //384pi/512
   m_sin[385]  =  11'b11001110000;     //385pi/512
   m_cos[385]  =  11'b11011000001;     //385pi/512
   m_sin[386]  =  11'b11001110010;     //386pi/512
   m_cos[386]  =  11'b11010111110;     //386pi/512
   m_sin[387]  =  11'b11001110100;     //387pi/512
   m_cos[387]  =  11'b11010111100;     //387pi/512
   m_sin[388]  =  11'b11001110101;     //388pi/512
   m_cos[388]  =  11'b11010111010;     //388pi/512
   m_sin[389]  =  11'b11001110111;     //389pi/512
   m_cos[389]  =  11'b11010110111;     //389pi/512
   m_sin[390]  =  11'b11001111001;     //390pi/512
   m_cos[390]  =  11'b11010110101;     //390pi/512
   m_sin[391]  =  11'b11001111011;     //391pi/512
   m_cos[391]  =  11'b11010110011;     //391pi/512
   m_sin[392]  =  11'b11001111101;     //392pi/512
   m_cos[392]  =  11'b11010110001;     //392pi/512
   m_sin[393]  =  11'b11001111111;     //393pi/512
   m_cos[393]  =  11'b11010101110;     //393pi/512
   m_sin[394]  =  11'b11010000001;     //394pi/512
   m_cos[394]  =  11'b11010101100;     //394pi/512
   m_sin[395]  =  11'b11010000011;     //395pi/512
   m_cos[395]  =  11'b11010101010;     //395pi/512
   m_sin[396]  =  11'b11010000101;     //396pi/512
   m_cos[396]  =  11'b11010101000;     //396pi/512
   m_sin[397]  =  11'b11010000111;     //397pi/512
   m_cos[397]  =  11'b11010100101;     //397pi/512
   m_sin[398]  =  11'b11010001001;     //398pi/512
   m_cos[398]  =  11'b11010100011;     //398pi/512
   m_sin[399]  =  11'b11010001011;     //399pi/512
   m_cos[399]  =  11'b11010100001;     //399pi/512
   m_sin[400]  =  11'b11010001101;     //400pi/512
   m_cos[400]  =  11'b11010011111;     //400pi/512
   m_sin[401]  =  11'b11010001111;     //401pi/512
   m_cos[401]  =  11'b11010011101;     //401pi/512
   m_sin[402]  =  11'b11010010001;     //402pi/512
   m_cos[402]  =  11'b11010011011;     //402pi/512
   m_sin[403]  =  11'b11010010011;     //403pi/512
   m_cos[403]  =  11'b11010011001;     //403pi/512
   m_sin[404]  =  11'b11010010110;     //404pi/512
   m_cos[404]  =  11'b11010010110;     //404pi/512
   m_sin[405]  =  11'b11010011000;     //405pi/512
   m_cos[405]  =  11'b11010010100;     //405pi/512
   m_sin[406]  =  11'b11010011010;     //406pi/512
   m_cos[406]  =  11'b11010010010;     //406pi/512
   m_sin[407]  =  11'b11010011100;     //407pi/512
   m_cos[407]  =  11'b11010010000;     //407pi/512
   m_sin[408]  =  11'b11010011110;     //408pi/512
   m_cos[408]  =  11'b11010001110;     //408pi/512
   m_sin[409]  =  11'b11010100000;     //409pi/512
   m_cos[409]  =  11'b11010001100;     //409pi/512
   m_sin[410]  =  11'b11010100010;     //410pi/512
   m_cos[410]  =  11'b11010001010;     //410pi/512
   m_sin[411]  =  11'b11010100101;     //411pi/512
   m_cos[411]  =  11'b11010001000;     //411pi/512
   m_sin[412]  =  11'b11010100111;     //412pi/512
   m_cos[412]  =  11'b11010000110;     //412pi/512
   m_sin[413]  =  11'b11010101001;     //413pi/512
   m_cos[413]  =  11'b11010000100;     //413pi/512
   m_sin[414]  =  11'b11010101011;     //414pi/512
   m_cos[414]  =  11'b11010000010;     //414pi/512
   m_sin[415]  =  11'b11010101101;     //415pi/512
   m_cos[415]  =  11'b11010000000;     //415pi/512
   m_sin[416]  =  11'b11010110000;     //416pi/512
   m_cos[416]  =  11'b11001111110;     //416pi/512
   m_sin[417]  =  11'b11010110010;     //417pi/512
   m_cos[417]  =  11'b11001111100;     //417pi/512
   m_sin[418]  =  11'b11010110100;     //418pi/512
   m_cos[418]  =  11'b11001111010;     //418pi/512
   m_sin[419]  =  11'b11010110110;     //419pi/512
   m_cos[419]  =  11'b11001111000;     //419pi/512
   m_sin[420]  =  11'b11010111001;     //420pi/512
   m_cos[420]  =  11'b11001110110;     //420pi/512
   m_sin[421]  =  11'b11010111011;     //421pi/512
   m_cos[421]  =  11'b11001110100;     //421pi/512
   m_sin[422]  =  11'b11010111101;     //422pi/512
   m_cos[422]  =  11'b11001110010;     //422pi/512
   m_sin[423]  =  11'b11011000000;     //423pi/512
   m_cos[423]  =  11'b11001110001;     //423pi/512
   m_sin[424]  =  11'b11011000010;     //424pi/512
   m_cos[424]  =  11'b11001101111;     //424pi/512
   m_sin[425]  =  11'b11011000100;     //425pi/512
   m_cos[425]  =  11'b11001101101;     //425pi/512
   m_sin[426]  =  11'b11011000111;     //426pi/512
   m_cos[426]  =  11'b11001101011;     //426pi/512
   m_sin[427]  =  11'b11011001001;     //427pi/512
   m_cos[427]  =  11'b11001101001;     //427pi/512
   m_sin[428]  =  11'b11011001011;     //428pi/512
   m_cos[428]  =  11'b11001100111;     //428pi/512
   m_sin[429]  =  11'b11011001110;     //429pi/512
   m_cos[429]  =  11'b11001100110;     //429pi/512
   m_sin[430]  =  11'b11011010000;     //430pi/512
   m_cos[430]  =  11'b11001100100;     //430pi/512
   m_sin[431]  =  11'b11011010011;     //431pi/512
   m_cos[431]  =  11'b11001100010;     //431pi/512
   m_sin[432]  =  11'b11011010101;     //432pi/512
   m_cos[432]  =  11'b11001100000;     //432pi/512
   m_sin[433]  =  11'b11011011000;     //433pi/512
   m_cos[433]  =  11'b11001011111;     //433pi/512
   m_sin[434]  =  11'b11011011010;     //434pi/512
   m_cos[434]  =  11'b11001011101;     //434pi/512
   m_sin[435]  =  11'b11011011100;     //435pi/512
   m_cos[435]  =  11'b11001011011;     //435pi/512
   m_sin[436]  =  11'b11011011111;     //436pi/512
   m_cos[436]  =  11'b11001011001;     //436pi/512
   m_sin[437]  =  11'b11011100001;     //437pi/512
   m_cos[437]  =  11'b11001011000;     //437pi/512
   m_sin[438]  =  11'b11011100100;     //438pi/512
   m_cos[438]  =  11'b11001010110;     //438pi/512
   m_sin[439]  =  11'b11011100110;     //439pi/512
   m_cos[439]  =  11'b11001010100;     //439pi/512
   m_sin[440]  =  11'b11011101001;     //440pi/512
   m_cos[440]  =  11'b11001010011;     //440pi/512
   m_sin[441]  =  11'b11011101011;     //441pi/512
   m_cos[441]  =  11'b11001010001;     //441pi/512
   m_sin[442]  =  11'b11011101110;     //442pi/512
   m_cos[442]  =  11'b11001010000;     //442pi/512
   m_sin[443]  =  11'b11011110000;     //443pi/512
   m_cos[443]  =  11'b11001001110;     //443pi/512
   m_sin[444]  =  11'b11011110011;     //444pi/512
   m_cos[444]  =  11'b11001001100;     //444pi/512
   m_sin[445]  =  11'b11011110101;     //445pi/512
   m_cos[445]  =  11'b11001001011;     //445pi/512
   m_sin[446]  =  11'b11011111000;     //446pi/512
   m_cos[446]  =  11'b11001001001;     //446pi/512
   m_sin[447]  =  11'b11011111011;     //447pi/512
   m_cos[447]  =  11'b11001001000;     //447pi/512
   m_sin[448]  =  11'b11011111101;     //448pi/512
   m_cos[448]  =  11'b11001000110;     //448pi/512
   m_sin[449]  =  11'b11100000000;     //449pi/512
   m_cos[449]  =  11'b11001000101;     //449pi/512
   m_sin[450]  =  11'b11100000010;     //450pi/512
   m_cos[450]  =  11'b11001000011;     //450pi/512
   m_sin[451]  =  11'b11100000101;     //451pi/512
   m_cos[451]  =  11'b11001000010;     //451pi/512
   m_sin[452]  =  11'b11100000111;     //452pi/512
   m_cos[452]  =  11'b11001000000;     //452pi/512
   m_sin[453]  =  11'b11100001010;     //453pi/512
   m_cos[453]  =  11'b11000111111;     //453pi/512
   m_sin[454]  =  11'b11100001101;     //454pi/512
   m_cos[454]  =  11'b11000111101;     //454pi/512
   m_sin[455]  =  11'b11100001111;     //455pi/512
   m_cos[455]  =  11'b11000111100;     //455pi/512
   m_sin[456]  =  11'b11100010010;     //456pi/512
   m_cos[456]  =  11'b11000111011;     //456pi/512
   m_sin[457]  =  11'b11100010101;     //457pi/512
   m_cos[457]  =  11'b11000111001;     //457pi/512
   m_sin[458]  =  11'b11100010111;     //458pi/512
   m_cos[458]  =  11'b11000111000;     //458pi/512
   m_sin[459]  =  11'b11100011010;     //459pi/512
   m_cos[459]  =  11'b11000110111;     //459pi/512
   m_sin[460]  =  11'b11100011101;     //460pi/512
   m_cos[460]  =  11'b11000110101;     //460pi/512
   m_sin[461]  =  11'b11100011111;     //461pi/512
   m_cos[461]  =  11'b11000110100;     //461pi/512
   m_sin[462]  =  11'b11100100010;     //462pi/512
   m_cos[462]  =  11'b11000110011;     //462pi/512
   m_sin[463]  =  11'b11100100101;     //463pi/512
   m_cos[463]  =  11'b11000110001;     //463pi/512
   m_sin[464]  =  11'b11100100111;     //464pi/512
   m_cos[464]  =  11'b11000110000;     //464pi/512
   m_sin[465]  =  11'b11100101010;     //465pi/512
   m_cos[465]  =  11'b11000101111;     //465pi/512
   m_sin[466]  =  11'b11100101101;     //466pi/512
   m_cos[466]  =  11'b11000101110;     //466pi/512
   m_sin[467]  =  11'b11100110000;     //467pi/512
   m_cos[467]  =  11'b11000101100;     //467pi/512
   m_sin[468]  =  11'b11100110010;     //468pi/512
   m_cos[468]  =  11'b11000101011;     //468pi/512
   m_sin[469]  =  11'b11100110101;     //469pi/512
   m_cos[469]  =  11'b11000101010;     //469pi/512
   m_sin[470]  =  11'b11100111000;     //470pi/512
   m_cos[470]  =  11'b11000101001;     //470pi/512
   m_sin[471]  =  11'b11100111010;     //471pi/512
   m_cos[471]  =  11'b11000101000;     //471pi/512
   m_sin[472]  =  11'b11100111101;     //472pi/512
   m_cos[472]  =  11'b11000100110;     //472pi/512
   m_sin[473]  =  11'b11101000000;     //473pi/512
   m_cos[473]  =  11'b11000100101;     //473pi/512
   m_sin[474]  =  11'b11101000011;     //474pi/512
   m_cos[474]  =  11'b11000100100;     //474pi/512
   m_sin[475]  =  11'b11101000110;     //475pi/512
   m_cos[475]  =  11'b11000100011;     //475pi/512
   m_sin[476]  =  11'b11101001000;     //476pi/512
   m_cos[476]  =  11'b11000100010;     //476pi/512
   m_sin[477]  =  11'b11101001011;     //477pi/512
   m_cos[477]  =  11'b11000100001;     //477pi/512
   m_sin[478]  =  11'b11101001110;     //478pi/512
   m_cos[478]  =  11'b11000100000;     //478pi/512
   m_sin[479]  =  11'b11101010001;     //479pi/512
   m_cos[479]  =  11'b11000011111;     //479pi/512
   m_sin[480]  =  11'b11101010100;     //480pi/512
   m_cos[480]  =  11'b11000011110;     //480pi/512
   m_sin[481]  =  11'b11101010110;     //481pi/512
   m_cos[481]  =  11'b11000011101;     //481pi/512
   m_sin[482]  =  11'b11101011001;     //482pi/512
   m_cos[482]  =  11'b11000011100;     //482pi/512
   m_sin[483]  =  11'b11101011100;     //483pi/512
   m_cos[483]  =  11'b11000011011;     //483pi/512
   m_sin[484]  =  11'b11101011111;     //484pi/512
   m_cos[484]  =  11'b11000011010;     //484pi/512
   m_sin[485]  =  11'b11101100010;     //485pi/512
   m_cos[485]  =  11'b11000011001;     //485pi/512
   m_sin[486]  =  11'b11101100100;     //486pi/512
   m_cos[486]  =  11'b11000011000;     //486pi/512
   m_sin[487]  =  11'b11101100111;     //487pi/512
   m_cos[487]  =  11'b11000010111;     //487pi/512
   m_sin[488]  =  11'b11101101010;     //488pi/512
   m_cos[488]  =  11'b11000010110;     //488pi/512
   m_sin[489]  =  11'b11101101101;     //489pi/512
   m_cos[489]  =  11'b11000010110;     //489pi/512
   m_sin[490]  =  11'b11101110000;     //490pi/512
   m_cos[490]  =  11'b11000010101;     //490pi/512
   m_sin[491]  =  11'b11101110011;     //491pi/512
   m_cos[491]  =  11'b11000010100;     //491pi/512
   m_sin[492]  =  11'b11101110110;     //492pi/512
   m_cos[492]  =  11'b11000010011;     //492pi/512
   m_sin[493]  =  11'b11101111001;     //493pi/512
   m_cos[493]  =  11'b11000010010;     //493pi/512
   m_sin[494]  =  11'b11101111011;     //494pi/512
   m_cos[494]  =  11'b11000010001;     //494pi/512
   m_sin[495]  =  11'b11101111110;     //495pi/512
   m_cos[495]  =  11'b11000010001;     //495pi/512
   m_sin[496]  =  11'b11110000001;     //496pi/512
   m_cos[496]  =  11'b11000010000;     //496pi/512
   m_sin[497]  =  11'b11110000100;     //497pi/512
   m_cos[497]  =  11'b11000001111;     //497pi/512
   m_sin[498]  =  11'b11110000111;     //498pi/512
   m_cos[498]  =  11'b11000001111;     //498pi/512
   m_sin[499]  =  11'b11110001010;     //499pi/512
   m_cos[499]  =  11'b11000001110;     //499pi/512
   m_sin[500]  =  11'b11110001101;     //500pi/512
   m_cos[500]  =  11'b11000001101;     //500pi/512
   m_sin[501]  =  11'b11110010000;     //501pi/512
   m_cos[501]  =  11'b11000001100;     //501pi/512
   m_sin[502]  =  11'b11110010011;     //502pi/512
   m_cos[502]  =  11'b11000001100;     //502pi/512
   m_sin[503]  =  11'b11110010101;     //503pi/512
   m_cos[503]  =  11'b11000001011;     //503pi/512
   m_sin[504]  =  11'b11110011000;     //504pi/512
   m_cos[504]  =  11'b11000001011;     //504pi/512
   m_sin[505]  =  11'b11110011011;     //505pi/512
   m_cos[505]  =  11'b11000001010;     //505pi/512
   m_sin[506]  =  11'b11110011110;     //506pi/512
   m_cos[506]  =  11'b11000001001;     //506pi/512
   m_sin[507]  =  11'b11110100001;     //507pi/512
   m_cos[507]  =  11'b11000001001;     //507pi/512
   m_sin[508]  =  11'b11110100100;     //508pi/512
   m_cos[508]  =  11'b11000001000;     //508pi/512
   m_sin[509]  =  11'b11110100111;     //509pi/512
   m_cos[509]  =  11'b11000001000;     //509pi/512
   m_sin[510]  =  11'b11110101010;     //510pi/512
   m_cos[510]  =  11'b11000000111;     //510pi/512
   m_sin[511]  =  11'b11110101101;     //511pi/512
   m_cos[511]  =  11'b11000000111;     //511pi/512
end
endmodule
