module  TWIDLE_10_bit  (
    input   [10:0]   rd_ptr_angle,

    output  signed [9:0]   cos_data,
    output  signed [9:0]   sin_data
 );

wire signed [9:0]  cos  [511:0];
wire signed [9:0]  sin  [511:0];

assign cos_data =    cos [rd_ptr_angle];
assign sin_data =    sin [rd_ptr_angle];

  assign sin[0]  =  10'b0000000000;     //0pi/512
  assign cos[0]  =  10'b0100000000;     //0pi/512
  assign sin[1]  =  10'b1111111110;     //1pi/512
  assign cos[1]  =  10'b0011111111;     //1pi/512
  assign sin[2]  =  10'b1111111101;     //2pi/512
  assign cos[2]  =  10'b0011111111;     //2pi/512
  assign sin[3]  =  10'b1111111011;     //3pi/512
  assign cos[3]  =  10'b0011111111;     //3pi/512
  assign sin[4]  =  10'b1111111010;     //4pi/512
  assign cos[4]  =  10'b0011111111;     //4pi/512
  assign sin[5]  =  10'b1111111000;     //5pi/512
  assign cos[5]  =  10'b0011111111;     //5pi/512
  assign sin[6]  =  10'b1111110111;     //6pi/512
  assign cos[6]  =  10'b0011111111;     //6pi/512
  assign sin[7]  =  10'b1111110101;     //7pi/512
  assign cos[7]  =  10'b0011111111;     //7pi/512
  assign sin[8]  =  10'b1111110011;     //8pi/512
  assign cos[8]  =  10'b0011111111;     //8pi/512
  assign sin[9]  =  10'b1111110010;     //9pi/512
  assign cos[9]  =  10'b0011111111;     //9pi/512
  assign sin[10]  =  10'b1111110000;     //10pi/512
  assign cos[10]  =  10'b0011111111;     //10pi/512
  assign sin[11]  =  10'b1111101111;     //11pi/512
  assign cos[11]  =  10'b0011111111;     //11pi/512
  assign sin[12]  =  10'b1111101101;     //12pi/512
  assign cos[12]  =  10'b0011111111;     //12pi/512
  assign sin[13]  =  10'b1111101100;     //13pi/512
  assign cos[13]  =  10'b0011111111;     //13pi/512
  assign sin[14]  =  10'b1111101010;     //14pi/512
  assign cos[14]  =  10'b0011111111;     //14pi/512
  assign sin[15]  =  10'b1111101000;     //15pi/512
  assign cos[15]  =  10'b0011111110;     //15pi/512
  assign sin[16]  =  10'b1111100111;     //16pi/512
  assign cos[16]  =  10'b0011111110;     //16pi/512
  assign sin[17]  =  10'b1111100101;     //17pi/512
  assign cos[17]  =  10'b0011111110;     //17pi/512
  assign sin[18]  =  10'b1111100100;     //18pi/512
  assign cos[18]  =  10'b0011111110;     //18pi/512
  assign sin[19]  =  10'b1111100010;     //19pi/512
  assign cos[19]  =  10'b0011111110;     //19pi/512
  assign sin[20]  =  10'b1111100001;     //20pi/512
  assign cos[20]  =  10'b0011111110;     //20pi/512
  assign sin[21]  =  10'b1111011111;     //21pi/512
  assign cos[21]  =  10'b0011111101;     //21pi/512
  assign sin[22]  =  10'b1111011110;     //22pi/512
  assign cos[22]  =  10'b0011111101;     //22pi/512
  assign sin[23]  =  10'b1111011100;     //23pi/512
  assign cos[23]  =  10'b0011111101;     //23pi/512
  assign sin[24]  =  10'b1111011010;     //24pi/512
  assign cos[24]  =  10'b0011111101;     //24pi/512
  assign sin[25]  =  10'b1111011001;     //25pi/512
  assign cos[25]  =  10'b0011111100;     //25pi/512
  assign sin[26]  =  10'b1111010111;     //26pi/512
  assign cos[26]  =  10'b0011111100;     //26pi/512
  assign sin[27]  =  10'b1111010110;     //27pi/512
  assign cos[27]  =  10'b0011111100;     //27pi/512
  assign sin[28]  =  10'b1111010100;     //28pi/512
  assign cos[28]  =  10'b0011111100;     //28pi/512
  assign sin[29]  =  10'b1111010011;     //29pi/512
  assign cos[29]  =  10'b0011111011;     //29pi/512
  assign sin[30]  =  10'b1111010001;     //30pi/512
  assign cos[30]  =  10'b0011111011;     //30pi/512
  assign sin[31]  =  10'b1111010000;     //31pi/512
  assign cos[31]  =  10'b0011111011;     //31pi/512
  assign sin[32]  =  10'b1111001110;     //32pi/512
  assign cos[32]  =  10'b0011111011;     //32pi/512
  assign sin[33]  =  10'b1111001101;     //33pi/512
  assign cos[33]  =  10'b0011111010;     //33pi/512
  assign sin[34]  =  10'b1111001011;     //34pi/512
  assign cos[34]  =  10'b0011111010;     //34pi/512
  assign sin[35]  =  10'b1111001001;     //35pi/512
  assign cos[35]  =  10'b0011111010;     //35pi/512
  assign sin[36]  =  10'b1111001000;     //36pi/512
  assign cos[36]  =  10'b0011111001;     //36pi/512
  assign sin[37]  =  10'b1111000110;     //37pi/512
  assign cos[37]  =  10'b0011111001;     //37pi/512
  assign sin[38]  =  10'b1111000101;     //38pi/512
  assign cos[38]  =  10'b0011111001;     //38pi/512
  assign sin[39]  =  10'b1111000011;     //39pi/512
  assign cos[39]  =  10'b0011111000;     //39pi/512
  assign sin[40]  =  10'b1111000010;     //40pi/512
  assign cos[40]  =  10'b0011111000;     //40pi/512
  assign sin[41]  =  10'b1111000000;     //41pi/512
  assign cos[41]  =  10'b0011110111;     //41pi/512
  assign sin[42]  =  10'b1110111111;     //42pi/512
  assign cos[42]  =  10'b0011110111;     //42pi/512
  assign sin[43]  =  10'b1110111101;     //43pi/512
  assign cos[43]  =  10'b0011110111;     //43pi/512
  assign sin[44]  =  10'b1110111100;     //44pi/512
  assign cos[44]  =  10'b0011110110;     //44pi/512
  assign sin[45]  =  10'b1110111010;     //45pi/512
  assign cos[45]  =  10'b0011110110;     //45pi/512
  assign sin[46]  =  10'b1110111001;     //46pi/512
  assign cos[46]  =  10'b0011110101;     //46pi/512
  assign sin[47]  =  10'b1110110111;     //47pi/512
  assign cos[47]  =  10'b0011110101;     //47pi/512
  assign sin[48]  =  10'b1110110110;     //48pi/512
  assign cos[48]  =  10'b0011110100;     //48pi/512
  assign sin[49]  =  10'b1110110100;     //49pi/512
  assign cos[49]  =  10'b0011110100;     //49pi/512
  assign sin[50]  =  10'b1110110011;     //50pi/512
  assign cos[50]  =  10'b0011110100;     //50pi/512
  assign sin[51]  =  10'b1110110001;     //51pi/512
  assign cos[51]  =  10'b0011110011;     //51pi/512
  assign sin[52]  =  10'b1110110000;     //52pi/512
  assign cos[52]  =  10'b0011110011;     //52pi/512
  assign sin[53]  =  10'b1110101110;     //53pi/512
  assign cos[53]  =  10'b0011110010;     //53pi/512
  assign sin[54]  =  10'b1110101101;     //54pi/512
  assign cos[54]  =  10'b0011110010;     //54pi/512
  assign sin[55]  =  10'b1110101011;     //55pi/512
  assign cos[55]  =  10'b0011110001;     //55pi/512
  assign sin[56]  =  10'b1110101010;     //56pi/512
  assign cos[56]  =  10'b0011110001;     //56pi/512
  assign sin[57]  =  10'b1110101000;     //57pi/512
  assign cos[57]  =  10'b0011110000;     //57pi/512
  assign sin[58]  =  10'b1110100111;     //58pi/512
  assign cos[58]  =  10'b0011101111;     //58pi/512
  assign sin[59]  =  10'b1110100101;     //59pi/512
  assign cos[59]  =  10'b0011101111;     //59pi/512
  assign sin[60]  =  10'b1110100100;     //60pi/512
  assign cos[60]  =  10'b0011101110;     //60pi/512
  assign sin[61]  =  10'b1110100010;     //61pi/512
  assign cos[61]  =  10'b0011101110;     //61pi/512
  assign sin[62]  =  10'b1110100001;     //62pi/512
  assign cos[62]  =  10'b0011101101;     //62pi/512
  assign sin[63]  =  10'b1110011111;     //63pi/512
  assign cos[63]  =  10'b0011101101;     //63pi/512
  assign sin[64]  =  10'b1110011110;     //64pi/512
  assign cos[64]  =  10'b0011101100;     //64pi/512
  assign sin[65]  =  10'b1110011101;     //65pi/512
  assign cos[65]  =  10'b0011101011;     //65pi/512
  assign sin[66]  =  10'b1110011011;     //66pi/512
  assign cos[66]  =  10'b0011101011;     //66pi/512
  assign sin[67]  =  10'b1110011010;     //67pi/512
  assign cos[67]  =  10'b0011101010;     //67pi/512
  assign sin[68]  =  10'b1110011000;     //68pi/512
  assign cos[68]  =  10'b0011101010;     //68pi/512
  assign sin[69]  =  10'b1110010111;     //69pi/512
  assign cos[69]  =  10'b0011101001;     //69pi/512
  assign sin[70]  =  10'b1110010101;     //70pi/512
  assign cos[70]  =  10'b0011101000;     //70pi/512
  assign sin[71]  =  10'b1110010100;     //71pi/512
  assign cos[71]  =  10'b0011101000;     //71pi/512
  assign sin[72]  =  10'b1110010011;     //72pi/512
  assign cos[72]  =  10'b0011100111;     //72pi/512
  assign sin[73]  =  10'b1110010001;     //73pi/512
  assign cos[73]  =  10'b0011100110;     //73pi/512
  assign sin[74]  =  10'b1110010000;     //74pi/512
  assign cos[74]  =  10'b0011100110;     //74pi/512
  assign sin[75]  =  10'b1110001110;     //75pi/512
  assign cos[75]  =  10'b0011100101;     //75pi/512
  assign sin[76]  =  10'b1110001101;     //76pi/512
  assign cos[76]  =  10'b0011100100;     //76pi/512
  assign sin[77]  =  10'b1110001011;     //77pi/512
  assign cos[77]  =  10'b0011100011;     //77pi/512
  assign sin[78]  =  10'b1110001010;     //78pi/512
  assign cos[78]  =  10'b0011100011;     //78pi/512
  assign sin[79]  =  10'b1110001001;     //79pi/512
  assign cos[79]  =  10'b0011100010;     //79pi/512
  assign sin[80]  =  10'b1110000111;     //80pi/512
  assign cos[80]  =  10'b0011100001;     //80pi/512
  assign sin[81]  =  10'b1110000110;     //81pi/512
  assign cos[81]  =  10'b0011100001;     //81pi/512
  assign sin[82]  =  10'b1110000101;     //82pi/512
  assign cos[82]  =  10'b0011100000;     //82pi/512
  assign sin[83]  =  10'b1110000011;     //83pi/512
  assign cos[83]  =  10'b0011011111;     //83pi/512
  assign sin[84]  =  10'b1110000010;     //84pi/512
  assign cos[84]  =  10'b0011011110;     //84pi/512
  assign sin[85]  =  10'b1110000000;     //85pi/512
  assign cos[85]  =  10'b0011011101;     //85pi/512
  assign sin[86]  =  10'b1101111111;     //86pi/512
  assign cos[86]  =  10'b0011011101;     //86pi/512
  assign sin[87]  =  10'b1101111110;     //87pi/512
  assign cos[87]  =  10'b0011011100;     //87pi/512
  assign sin[88]  =  10'b1101111100;     //88pi/512
  assign cos[88]  =  10'b0011011011;     //88pi/512
  assign sin[89]  =  10'b1101111011;     //89pi/512
  assign cos[89]  =  10'b0011011010;     //89pi/512
  assign sin[90]  =  10'b1101111010;     //90pi/512
  assign cos[90]  =  10'b0011011001;     //90pi/512
  assign sin[91]  =  10'b1101111000;     //91pi/512
  assign cos[91]  =  10'b0011011001;     //91pi/512
  assign sin[92]  =  10'b1101110111;     //92pi/512
  assign cos[92]  =  10'b0011011000;     //92pi/512
  assign sin[93]  =  10'b1101110110;     //93pi/512
  assign cos[93]  =  10'b0011010111;     //93pi/512
  assign sin[94]  =  10'b1101110100;     //94pi/512
  assign cos[94]  =  10'b0011010110;     //94pi/512
  assign sin[95]  =  10'b1101110011;     //95pi/512
  assign cos[95]  =  10'b0011010101;     //95pi/512
  assign sin[96]  =  10'b1101110010;     //96pi/512
  assign cos[96]  =  10'b0011010100;     //96pi/512
  assign sin[97]  =  10'b1101110000;     //97pi/512
  assign cos[97]  =  10'b0011010011;     //97pi/512
  assign sin[98]  =  10'b1101101111;     //98pi/512
  assign cos[98]  =  10'b0011010011;     //98pi/512
  assign sin[99]  =  10'b1101101110;     //99pi/512
  assign cos[99]  =  10'b0011010010;     //99pi/512
  assign sin[100]  =  10'b1101101101;     //100pi/512
  assign cos[100]  =  10'b0011010001;     //100pi/512
  assign sin[101]  =  10'b1101101011;     //101pi/512
  assign cos[101]  =  10'b0011010000;     //101pi/512
  assign sin[102]  =  10'b1101101010;     //102pi/512
  assign cos[102]  =  10'b0011001111;     //102pi/512
  assign sin[103]  =  10'b1101101001;     //103pi/512
  assign cos[103]  =  10'b0011001110;     //103pi/512
  assign sin[104]  =  10'b1101101000;     //104pi/512
  assign cos[104]  =  10'b0011001101;     //104pi/512
  assign sin[105]  =  10'b1101100110;     //105pi/512
  assign cos[105]  =  10'b0011001100;     //105pi/512
  assign sin[106]  =  10'b1101100101;     //106pi/512
  assign cos[106]  =  10'b0011001011;     //106pi/512
  assign sin[107]  =  10'b1101100100;     //107pi/512
  assign cos[107]  =  10'b0011001010;     //107pi/512
  assign sin[108]  =  10'b1101100011;     //108pi/512
  assign cos[108]  =  10'b0011001001;     //108pi/512
  assign sin[109]  =  10'b1101100001;     //109pi/512
  assign cos[109]  =  10'b0011001000;     //109pi/512
  assign sin[110]  =  10'b1101100000;     //110pi/512
  assign cos[110]  =  10'b0011000111;     //110pi/512
  assign sin[111]  =  10'b1101011111;     //111pi/512
  assign cos[111]  =  10'b0011000110;     //111pi/512
  assign sin[112]  =  10'b1101011110;     //112pi/512
  assign cos[112]  =  10'b0011000101;     //112pi/512
  assign sin[113]  =  10'b1101011100;     //113pi/512
  assign cos[113]  =  10'b0011000100;     //113pi/512
  assign sin[114]  =  10'b1101011011;     //114pi/512
  assign cos[114]  =  10'b0011000011;     //114pi/512
  assign sin[115]  =  10'b1101011010;     //115pi/512
  assign cos[115]  =  10'b0011000010;     //115pi/512
  assign sin[116]  =  10'b1101011001;     //116pi/512
  assign cos[116]  =  10'b0011000001;     //116pi/512
  assign sin[117]  =  10'b1101011000;     //117pi/512
  assign cos[117]  =  10'b0011000000;     //117pi/512
  assign sin[118]  =  10'b1101010110;     //118pi/512
  assign cos[118]  =  10'b0010111111;     //118pi/512
  assign sin[119]  =  10'b1101010101;     //119pi/512
  assign cos[119]  =  10'b0010111110;     //119pi/512
  assign sin[120]  =  10'b1101010100;     //120pi/512
  assign cos[120]  =  10'b0010111101;     //120pi/512
  assign sin[121]  =  10'b1101010011;     //121pi/512
  assign cos[121]  =  10'b0010111100;     //121pi/512
  assign sin[122]  =  10'b1101010010;     //122pi/512
  assign cos[122]  =  10'b0010111011;     //122pi/512
  assign sin[123]  =  10'b1101010001;     //123pi/512
  assign cos[123]  =  10'b0010111010;     //123pi/512
  assign sin[124]  =  10'b1101001111;     //124pi/512
  assign cos[124]  =  10'b0010111001;     //124pi/512
  assign sin[125]  =  10'b1101001110;     //125pi/512
  assign cos[125]  =  10'b0010111000;     //125pi/512
  assign sin[126]  =  10'b1101001101;     //126pi/512
  assign cos[126]  =  10'b0010110111;     //126pi/512
  assign sin[127]  =  10'b1101001100;     //127pi/512
  assign cos[127]  =  10'b0010110110;     //127pi/512
  assign sin[128]  =  10'b1101001011;     //128pi/512
  assign cos[128]  =  10'b0010110101;     //128pi/512
  assign sin[129]  =  10'b1101001010;     //129pi/512
  assign cos[129]  =  10'b0010110011;     //129pi/512
  assign sin[130]  =  10'b1101001001;     //130pi/512
  assign cos[130]  =  10'b0010110010;     //130pi/512
  assign sin[131]  =  10'b1101001000;     //131pi/512
  assign cos[131]  =  10'b0010110001;     //131pi/512
  assign sin[132]  =  10'b1101000111;     //132pi/512
  assign cos[132]  =  10'b0010110000;     //132pi/512
  assign sin[133]  =  10'b1101000110;     //133pi/512
  assign cos[133]  =  10'b0010101111;     //133pi/512
  assign sin[134]  =  10'b1101000100;     //134pi/512
  assign cos[134]  =  10'b0010101110;     //134pi/512
  assign sin[135]  =  10'b1101000011;     //135pi/512
  assign cos[135]  =  10'b0010101101;     //135pi/512
  assign sin[136]  =  10'b1101000010;     //136pi/512
  assign cos[136]  =  10'b0010101011;     //136pi/512
  assign sin[137]  =  10'b1101000001;     //137pi/512
  assign cos[137]  =  10'b0010101010;     //137pi/512
  assign sin[138]  =  10'b1101000000;     //138pi/512
  assign cos[138]  =  10'b0010101001;     //138pi/512
  assign sin[139]  =  10'b1100111111;     //139pi/512
  assign cos[139]  =  10'b0010101000;     //139pi/512
  assign sin[140]  =  10'b1100111110;     //140pi/512
  assign cos[140]  =  10'b0010100111;     //140pi/512
  assign sin[141]  =  10'b1100111101;     //141pi/512
  assign cos[141]  =  10'b0010100110;     //141pi/512
  assign sin[142]  =  10'b1100111100;     //142pi/512
  assign cos[142]  =  10'b0010100100;     //142pi/512
  assign sin[143]  =  10'b1100111011;     //143pi/512
  assign cos[143]  =  10'b0010100011;     //143pi/512
  assign sin[144]  =  10'b1100111010;     //144pi/512
  assign cos[144]  =  10'b0010100010;     //144pi/512
  assign sin[145]  =  10'b1100111001;     //145pi/512
  assign cos[145]  =  10'b0010100001;     //145pi/512
  assign sin[146]  =  10'b1100111000;     //146pi/512
  assign cos[146]  =  10'b0010011111;     //146pi/512
  assign sin[147]  =  10'b1100110111;     //147pi/512
  assign cos[147]  =  10'b0010011110;     //147pi/512
  assign sin[148]  =  10'b1100110110;     //148pi/512
  assign cos[148]  =  10'b0010011101;     //148pi/512
  assign sin[149]  =  10'b1100110101;     //149pi/512
  assign cos[149]  =  10'b0010011100;     //149pi/512
  assign sin[150]  =  10'b1100110100;     //150pi/512
  assign cos[150]  =  10'b0010011011;     //150pi/512
  assign sin[151]  =  10'b1100110011;     //151pi/512
  assign cos[151]  =  10'b0010011001;     //151pi/512
  assign sin[152]  =  10'b1100110010;     //152pi/512
  assign cos[152]  =  10'b0010011000;     //152pi/512
  assign sin[153]  =  10'b1100110001;     //153pi/512
  assign cos[153]  =  10'b0010010111;     //153pi/512
  assign sin[154]  =  10'b1100110001;     //154pi/512
  assign cos[154]  =  10'b0010010101;     //154pi/512
  assign sin[155]  =  10'b1100110000;     //155pi/512
  assign cos[155]  =  10'b0010010100;     //155pi/512
  assign sin[156]  =  10'b1100101111;     //156pi/512
  assign cos[156]  =  10'b0010010011;     //156pi/512
  assign sin[157]  =  10'b1100101110;     //157pi/512
  assign cos[157]  =  10'b0010010010;     //157pi/512
  assign sin[158]  =  10'b1100101101;     //158pi/512
  assign cos[158]  =  10'b0010010000;     //158pi/512
  assign sin[159]  =  10'b1100101100;     //159pi/512
  assign cos[159]  =  10'b0010001111;     //159pi/512
  assign sin[160]  =  10'b1100101011;     //160pi/512
  assign cos[160]  =  10'b0010001110;     //160pi/512
  assign sin[161]  =  10'b1100101010;     //161pi/512
  assign cos[161]  =  10'b0010001100;     //161pi/512
  assign sin[162]  =  10'b1100101001;     //162pi/512
  assign cos[162]  =  10'b0010001011;     //162pi/512
  assign sin[163]  =  10'b1100101001;     //163pi/512
  assign cos[163]  =  10'b0010001010;     //163pi/512
  assign sin[164]  =  10'b1100101000;     //164pi/512
  assign cos[164]  =  10'b0010001000;     //164pi/512
  assign sin[165]  =  10'b1100100111;     //165pi/512
  assign cos[165]  =  10'b0010000111;     //165pi/512
  assign sin[166]  =  10'b1100100110;     //166pi/512
  assign cos[166]  =  10'b0010000110;     //166pi/512
  assign sin[167]  =  10'b1100100101;     //167pi/512
  assign cos[167]  =  10'b0010000100;     //167pi/512
  assign sin[168]  =  10'b1100100100;     //168pi/512
  assign cos[168]  =  10'b0010000011;     //168pi/512
  assign sin[169]  =  10'b1100100100;     //169pi/512
  assign cos[169]  =  10'b0010000010;     //169pi/512
  assign sin[170]  =  10'b1100100011;     //170pi/512
  assign cos[170]  =  10'b0010000000;     //170pi/512
  assign sin[171]  =  10'b1100100010;     //171pi/512
  assign cos[171]  =  10'b0001111111;     //171pi/512
  assign sin[172]  =  10'b1100100001;     //172pi/512
  assign cos[172]  =  10'b0001111110;     //172pi/512
  assign sin[173]  =  10'b1100100000;     //173pi/512
  assign cos[173]  =  10'b0001111100;     //173pi/512
  assign sin[174]  =  10'b1100100000;     //174pi/512
  assign cos[174]  =  10'b0001111011;     //174pi/512
  assign sin[175]  =  10'b1100011111;     //175pi/512
  assign cos[175]  =  10'b0001111010;     //175pi/512
  assign sin[176]  =  10'b1100011110;     //176pi/512
  assign cos[176]  =  10'b0001111000;     //176pi/512
  assign sin[177]  =  10'b1100011101;     //177pi/512
  assign cos[177]  =  10'b0001110111;     //177pi/512
  assign sin[178]  =  10'b1100011101;     //178pi/512
  assign cos[178]  =  10'b0001110101;     //178pi/512
  assign sin[179]  =  10'b1100011100;     //179pi/512
  assign cos[179]  =  10'b0001110100;     //179pi/512
  assign sin[180]  =  10'b1100011011;     //180pi/512
  assign cos[180]  =  10'b0001110011;     //180pi/512
  assign sin[181]  =  10'b1100011011;     //181pi/512
  assign cos[181]  =  10'b0001110001;     //181pi/512
  assign sin[182]  =  10'b1100011010;     //182pi/512
  assign cos[182]  =  10'b0001110000;     //182pi/512
  assign sin[183]  =  10'b1100011001;     //183pi/512
  assign cos[183]  =  10'b0001101110;     //183pi/512
  assign sin[184]  =  10'b1100011001;     //184pi/512
  assign cos[184]  =  10'b0001101101;     //184pi/512
  assign sin[185]  =  10'b1100011000;     //185pi/512
  assign cos[185]  =  10'b0001101100;     //185pi/512
  assign sin[186]  =  10'b1100010111;     //186pi/512
  assign cos[186]  =  10'b0001101010;     //186pi/512
  assign sin[187]  =  10'b1100010111;     //187pi/512
  assign cos[187]  =  10'b0001101001;     //187pi/512
  assign sin[188]  =  10'b1100010110;     //188pi/512
  assign cos[188]  =  10'b0001100111;     //188pi/512
  assign sin[189]  =  10'b1100010101;     //189pi/512
  assign cos[189]  =  10'b0001100110;     //189pi/512
  assign sin[190]  =  10'b1100010101;     //190pi/512
  assign cos[190]  =  10'b0001100100;     //190pi/512
  assign sin[191]  =  10'b1100010100;     //191pi/512
  assign cos[191]  =  10'b0001100011;     //191pi/512
  assign sin[192]  =  10'b1100010011;     //192pi/512
  assign cos[192]  =  10'b0001100001;     //192pi/512
  assign sin[193]  =  10'b1100010011;     //193pi/512
  assign cos[193]  =  10'b0001100000;     //193pi/512
  assign sin[194]  =  10'b1100010010;     //194pi/512
  assign cos[194]  =  10'b0001011111;     //194pi/512
  assign sin[195]  =  10'b1100010010;     //195pi/512
  assign cos[195]  =  10'b0001011101;     //195pi/512
  assign sin[196]  =  10'b1100010001;     //196pi/512
  assign cos[196]  =  10'b0001011100;     //196pi/512
  assign sin[197]  =  10'b1100010001;     //197pi/512
  assign cos[197]  =  10'b0001011010;     //197pi/512
  assign sin[198]  =  10'b1100010000;     //198pi/512
  assign cos[198]  =  10'b0001011001;     //198pi/512
  assign sin[199]  =  10'b1100001111;     //199pi/512
  assign cos[199]  =  10'b0001010111;     //199pi/512
  assign sin[200]  =  10'b1100001111;     //200pi/512
  assign cos[200]  =  10'b0001010110;     //200pi/512
  assign sin[201]  =  10'b1100001110;     //201pi/512
  assign cos[201]  =  10'b0001010100;     //201pi/512
  assign sin[202]  =  10'b1100001110;     //202pi/512
  assign cos[202]  =  10'b0001010011;     //202pi/512
  assign sin[203]  =  10'b1100001101;     //203pi/512
  assign cos[203]  =  10'b0001010001;     //203pi/512
  assign sin[204]  =  10'b1100001101;     //204pi/512
  assign cos[204]  =  10'b0001010000;     //204pi/512
  assign sin[205]  =  10'b1100001100;     //205pi/512
  assign cos[205]  =  10'b0001001110;     //205pi/512
  assign sin[206]  =  10'b1100001100;     //206pi/512
  assign cos[206]  =  10'b0001001101;     //206pi/512
  assign sin[207]  =  10'b1100001011;     //207pi/512
  assign cos[207]  =  10'b0001001011;     //207pi/512
  assign sin[208]  =  10'b1100001011;     //208pi/512
  assign cos[208]  =  10'b0001001010;     //208pi/512
  assign sin[209]  =  10'b1100001011;     //209pi/512
  assign cos[209]  =  10'b0001001000;     //209pi/512
  assign sin[210]  =  10'b1100001010;     //210pi/512
  assign cos[210]  =  10'b0001000111;     //210pi/512
  assign sin[211]  =  10'b1100001010;     //211pi/512
  assign cos[211]  =  10'b0001000101;     //211pi/512
  assign sin[212]  =  10'b1100001001;     //212pi/512
  assign cos[212]  =  10'b0001000100;     //212pi/512
  assign sin[213]  =  10'b1100001001;     //213pi/512
  assign cos[213]  =  10'b0001000010;     //213pi/512
  assign sin[214]  =  10'b1100001000;     //214pi/512
  assign cos[214]  =  10'b0001000001;     //214pi/512
  assign sin[215]  =  10'b1100001000;     //215pi/512
  assign cos[215]  =  10'b0000111111;     //215pi/512
  assign sin[216]  =  10'b1100001000;     //216pi/512
  assign cos[216]  =  10'b0000111110;     //216pi/512
  assign sin[217]  =  10'b1100000111;     //217pi/512
  assign cos[217]  =  10'b0000111100;     //217pi/512
  assign sin[218]  =  10'b1100000111;     //218pi/512
  assign cos[218]  =  10'b0000111011;     //218pi/512
  assign sin[219]  =  10'b1100000111;     //219pi/512
  assign cos[219]  =  10'b0000111001;     //219pi/512
  assign sin[220]  =  10'b1100000110;     //220pi/512
  assign cos[220]  =  10'b0000111000;     //220pi/512
  assign sin[221]  =  10'b1100000110;     //221pi/512
  assign cos[221]  =  10'b0000110110;     //221pi/512
  assign sin[222]  =  10'b1100000110;     //222pi/512
  assign cos[222]  =  10'b0000110101;     //222pi/512
  assign sin[223]  =  10'b1100000101;     //223pi/512
  assign cos[223]  =  10'b0000110011;     //223pi/512
  assign sin[224]  =  10'b1100000101;     //224pi/512
  assign cos[224]  =  10'b0000110001;     //224pi/512
  assign sin[225]  =  10'b1100000101;     //225pi/512
  assign cos[225]  =  10'b0000110000;     //225pi/512
  assign sin[226]  =  10'b1100000100;     //226pi/512
  assign cos[226]  =  10'b0000101110;     //226pi/512
  assign sin[227]  =  10'b1100000100;     //227pi/512
  assign cos[227]  =  10'b0000101101;     //227pi/512
  assign sin[228]  =  10'b1100000100;     //228pi/512
  assign cos[228]  =  10'b0000101011;     //228pi/512
  assign sin[229]  =  10'b1100000100;     //229pi/512
  assign cos[229]  =  10'b0000101010;     //229pi/512
  assign sin[230]  =  10'b1100000011;     //230pi/512
  assign cos[230]  =  10'b0000101000;     //230pi/512
  assign sin[231]  =  10'b1100000011;     //231pi/512
  assign cos[231]  =  10'b0000100111;     //231pi/512
  assign sin[232]  =  10'b1100000011;     //232pi/512
  assign cos[232]  =  10'b0000100101;     //232pi/512
  assign sin[233]  =  10'b1100000011;     //233pi/512
  assign cos[233]  =  10'b0000100100;     //233pi/512
  assign sin[234]  =  10'b1100000010;     //234pi/512
  assign cos[234]  =  10'b0000100010;     //234pi/512
  assign sin[235]  =  10'b1100000010;     //235pi/512
  assign cos[235]  =  10'b0000100000;     //235pi/512
  assign sin[236]  =  10'b1100000010;     //236pi/512
  assign cos[236]  =  10'b0000011111;     //236pi/512
  assign sin[237]  =  10'b1100000010;     //237pi/512
  assign cos[237]  =  10'b0000011101;     //237pi/512
  assign sin[238]  =  10'b1100000010;     //238pi/512
  assign cos[238]  =  10'b0000011100;     //238pi/512
  assign sin[239]  =  10'b1100000001;     //239pi/512
  assign cos[239]  =  10'b0000011010;     //239pi/512
  assign sin[240]  =  10'b1100000001;     //240pi/512
  assign cos[240]  =  10'b0000011001;     //240pi/512
  assign sin[241]  =  10'b1100000001;     //241pi/512
  assign cos[241]  =  10'b0000010111;     //241pi/512
  assign sin[242]  =  10'b1100000001;     //242pi/512
  assign cos[242]  =  10'b0000010101;     //242pi/512
  assign sin[243]  =  10'b1100000001;     //243pi/512
  assign cos[243]  =  10'b0000010100;     //243pi/512
  assign sin[244]  =  10'b1100000001;     //244pi/512
  assign cos[244]  =  10'b0000010010;     //244pi/512
  assign sin[245]  =  10'b1100000001;     //245pi/512
  assign cos[245]  =  10'b0000010001;     //245pi/512
  assign sin[246]  =  10'b1100000000;     //246pi/512
  assign cos[246]  =  10'b0000001111;     //246pi/512
  assign sin[247]  =  10'b1100000000;     //247pi/512
  assign cos[247]  =  10'b0000001110;     //247pi/512
  assign sin[248]  =  10'b1100000000;     //248pi/512
  assign cos[248]  =  10'b0000001100;     //248pi/512
  assign sin[249]  =  10'b1100000000;     //249pi/512
  assign cos[249]  =  10'b0000001010;     //249pi/512
  assign sin[250]  =  10'b1100000000;     //250pi/512
  assign cos[250]  =  10'b0000001001;     //250pi/512
  assign sin[251]  =  10'b1100000000;     //251pi/512
  assign cos[251]  =  10'b0000000111;     //251pi/512
  assign sin[252]  =  10'b1100000000;     //252pi/512
  assign cos[252]  =  10'b0000000110;     //252pi/512
  assign sin[253]  =  10'b1100000000;     //253pi/512
  assign cos[253]  =  10'b0000000100;     //253pi/512
  assign sin[254]  =  10'b1100000000;     //254pi/512
  assign cos[254]  =  10'b0000000011;     //254pi/512
  assign sin[255]  =  10'b1100000000;     //255pi/512
  assign cos[255]  =  10'b0000000001;     //255pi/512
  assign sin[256]  =  10'b1100000000;     //256pi/512
  assign cos[256]  =  10'b0000000000;     //256pi/512
  assign sin[257]  =  10'b1100000000;     //257pi/512
  assign cos[257]  =  10'b1111111110;     //257pi/512
  assign sin[258]  =  10'b1100000000;     //258pi/512
  assign cos[258]  =  10'b1111111101;     //258pi/512
  assign sin[259]  =  10'b1100000000;     //259pi/512
  assign cos[259]  =  10'b1111111011;     //259pi/512
  assign sin[260]  =  10'b1100000000;     //260pi/512
  assign cos[260]  =  10'b1111111010;     //260pi/512
  assign sin[261]  =  10'b1100000000;     //261pi/512
  assign cos[261]  =  10'b1111111000;     //261pi/512
  assign sin[262]  =  10'b1100000000;     //262pi/512
  assign cos[262]  =  10'b1111110111;     //262pi/512
  assign sin[263]  =  10'b1100000000;     //263pi/512
  assign cos[263]  =  10'b1111110101;     //263pi/512
  assign sin[264]  =  10'b1100000000;     //264pi/512
  assign cos[264]  =  10'b1111110011;     //264pi/512
  assign sin[265]  =  10'b1100000000;     //265pi/512
  assign cos[265]  =  10'b1111110010;     //265pi/512
  assign sin[266]  =  10'b1100000000;     //266pi/512
  assign cos[266]  =  10'b1111110000;     //266pi/512
  assign sin[267]  =  10'b1100000001;     //267pi/512
  assign cos[267]  =  10'b1111101111;     //267pi/512
  assign sin[268]  =  10'b1100000001;     //268pi/512
  assign cos[268]  =  10'b1111101101;     //268pi/512
  assign sin[269]  =  10'b1100000001;     //269pi/512
  assign cos[269]  =  10'b1111101100;     //269pi/512
  assign sin[270]  =  10'b1100000001;     //270pi/512
  assign cos[270]  =  10'b1111101010;     //270pi/512
  assign sin[271]  =  10'b1100000001;     //271pi/512
  assign cos[271]  =  10'b1111101000;     //271pi/512
  assign sin[272]  =  10'b1100000001;     //272pi/512
  assign cos[272]  =  10'b1111100111;     //272pi/512
  assign sin[273]  =  10'b1100000001;     //273pi/512
  assign cos[273]  =  10'b1111100101;     //273pi/512
  assign sin[274]  =  10'b1100000010;     //274pi/512
  assign cos[274]  =  10'b1111100100;     //274pi/512
  assign sin[275]  =  10'b1100000010;     //275pi/512
  assign cos[275]  =  10'b1111100010;     //275pi/512
  assign sin[276]  =  10'b1100000010;     //276pi/512
  assign cos[276]  =  10'b1111100001;     //276pi/512
  assign sin[277]  =  10'b1100000010;     //277pi/512
  assign cos[277]  =  10'b1111011111;     //277pi/512
  assign sin[278]  =  10'b1100000010;     //278pi/512
  assign cos[278]  =  10'b1111011110;     //278pi/512
  assign sin[279]  =  10'b1100000011;     //279pi/512
  assign cos[279]  =  10'b1111011100;     //279pi/512
  assign sin[280]  =  10'b1100000011;     //280pi/512
  assign cos[280]  =  10'b1111011010;     //280pi/512
  assign sin[281]  =  10'b1100000011;     //281pi/512
  assign cos[281]  =  10'b1111011001;     //281pi/512
  assign sin[282]  =  10'b1100000011;     //282pi/512
  assign cos[282]  =  10'b1111010111;     //282pi/512
  assign sin[283]  =  10'b1100000100;     //283pi/512
  assign cos[283]  =  10'b1111010110;     //283pi/512
  assign sin[284]  =  10'b1100000100;     //284pi/512
  assign cos[284]  =  10'b1111010100;     //284pi/512
  assign sin[285]  =  10'b1100000100;     //285pi/512
  assign cos[285]  =  10'b1111010011;     //285pi/512
  assign sin[286]  =  10'b1100000100;     //286pi/512
  assign cos[286]  =  10'b1111010001;     //286pi/512
  assign sin[287]  =  10'b1100000101;     //287pi/512
  assign cos[287]  =  10'b1111010000;     //287pi/512
  assign sin[288]  =  10'b1100000101;     //288pi/512
  assign cos[288]  =  10'b1111001110;     //288pi/512
  assign sin[289]  =  10'b1100000101;     //289pi/512
  assign cos[289]  =  10'b1111001101;     //289pi/512
  assign sin[290]  =  10'b1100000110;     //290pi/512
  assign cos[290]  =  10'b1111001011;     //290pi/512
  assign sin[291]  =  10'b1100000110;     //291pi/512
  assign cos[291]  =  10'b1111001001;     //291pi/512
  assign sin[292]  =  10'b1100000110;     //292pi/512
  assign cos[292]  =  10'b1111001000;     //292pi/512
  assign sin[293]  =  10'b1100000111;     //293pi/512
  assign cos[293]  =  10'b1111000110;     //293pi/512
  assign sin[294]  =  10'b1100000111;     //294pi/512
  assign cos[294]  =  10'b1111000101;     //294pi/512
  assign sin[295]  =  10'b1100000111;     //295pi/512
  assign cos[295]  =  10'b1111000011;     //295pi/512
  assign sin[296]  =  10'b1100001000;     //296pi/512
  assign cos[296]  =  10'b1111000010;     //296pi/512
  assign sin[297]  =  10'b1100001000;     //297pi/512
  assign cos[297]  =  10'b1111000000;     //297pi/512
  assign sin[298]  =  10'b1100001000;     //298pi/512
  assign cos[298]  =  10'b1110111111;     //298pi/512
  assign sin[299]  =  10'b1100001001;     //299pi/512
  assign cos[299]  =  10'b1110111101;     //299pi/512
  assign sin[300]  =  10'b1100001001;     //300pi/512
  assign cos[300]  =  10'b1110111100;     //300pi/512
  assign sin[301]  =  10'b1100001010;     //301pi/512
  assign cos[301]  =  10'b1110111010;     //301pi/512
  assign sin[302]  =  10'b1100001010;     //302pi/512
  assign cos[302]  =  10'b1110111001;     //302pi/512
  assign sin[303]  =  10'b1100001011;     //303pi/512
  assign cos[303]  =  10'b1110110111;     //303pi/512
  assign sin[304]  =  10'b1100001011;     //304pi/512
  assign cos[304]  =  10'b1110110110;     //304pi/512
  assign sin[305]  =  10'b1100001011;     //305pi/512
  assign cos[305]  =  10'b1110110100;     //305pi/512
  assign sin[306]  =  10'b1100001100;     //306pi/512
  assign cos[306]  =  10'b1110110011;     //306pi/512
  assign sin[307]  =  10'b1100001100;     //307pi/512
  assign cos[307]  =  10'b1110110001;     //307pi/512
  assign sin[308]  =  10'b1100001101;     //308pi/512
  assign cos[308]  =  10'b1110110000;     //308pi/512
  assign sin[309]  =  10'b1100001101;     //309pi/512
  assign cos[309]  =  10'b1110101110;     //309pi/512
  assign sin[310]  =  10'b1100001110;     //310pi/512
  assign cos[310]  =  10'b1110101101;     //310pi/512
  assign sin[311]  =  10'b1100001110;     //311pi/512
  assign cos[311]  =  10'b1110101011;     //311pi/512
  assign sin[312]  =  10'b1100001111;     //312pi/512
  assign cos[312]  =  10'b1110101010;     //312pi/512
  assign sin[313]  =  10'b1100001111;     //313pi/512
  assign cos[313]  =  10'b1110101000;     //313pi/512
  assign sin[314]  =  10'b1100010000;     //314pi/512
  assign cos[314]  =  10'b1110100111;     //314pi/512
  assign sin[315]  =  10'b1100010001;     //315pi/512
  assign cos[315]  =  10'b1110100101;     //315pi/512
  assign sin[316]  =  10'b1100010001;     //316pi/512
  assign cos[316]  =  10'b1110100100;     //316pi/512
  assign sin[317]  =  10'b1100010010;     //317pi/512
  assign cos[317]  =  10'b1110100010;     //317pi/512
  assign sin[318]  =  10'b1100010010;     //318pi/512
  assign cos[318]  =  10'b1110100001;     //318pi/512
  assign sin[319]  =  10'b1100010011;     //319pi/512
  assign cos[319]  =  10'b1110011111;     //319pi/512
  assign sin[320]  =  10'b1100010011;     //320pi/512
  assign cos[320]  =  10'b1110011110;     //320pi/512
  assign sin[321]  =  10'b1100010100;     //321pi/512
  assign cos[321]  =  10'b1110011101;     //321pi/512
  assign sin[322]  =  10'b1100010101;     //322pi/512
  assign cos[322]  =  10'b1110011011;     //322pi/512
  assign sin[323]  =  10'b1100010101;     //323pi/512
  assign cos[323]  =  10'b1110011010;     //323pi/512
  assign sin[324]  =  10'b1100010110;     //324pi/512
  assign cos[324]  =  10'b1110011000;     //324pi/512
  assign sin[325]  =  10'b1100010111;     //325pi/512
  assign cos[325]  =  10'b1110010111;     //325pi/512
  assign sin[326]  =  10'b1100010111;     //326pi/512
  assign cos[326]  =  10'b1110010101;     //326pi/512
  assign sin[327]  =  10'b1100011000;     //327pi/512
  assign cos[327]  =  10'b1110010100;     //327pi/512
  assign sin[328]  =  10'b1100011001;     //328pi/512
  assign cos[328]  =  10'b1110010011;     //328pi/512
  assign sin[329]  =  10'b1100011001;     //329pi/512
  assign cos[329]  =  10'b1110010001;     //329pi/512
  assign sin[330]  =  10'b1100011010;     //330pi/512
  assign cos[330]  =  10'b1110010000;     //330pi/512
  assign sin[331]  =  10'b1100011011;     //331pi/512
  assign cos[331]  =  10'b1110001110;     //331pi/512
  assign sin[332]  =  10'b1100011011;     //332pi/512
  assign cos[332]  =  10'b1110001101;     //332pi/512
  assign sin[333]  =  10'b1100011100;     //333pi/512
  assign cos[333]  =  10'b1110001011;     //333pi/512
  assign sin[334]  =  10'b1100011101;     //334pi/512
  assign cos[334]  =  10'b1110001010;     //334pi/512
  assign sin[335]  =  10'b1100011101;     //335pi/512
  assign cos[335]  =  10'b1110001001;     //335pi/512
  assign sin[336]  =  10'b1100011110;     //336pi/512
  assign cos[336]  =  10'b1110000111;     //336pi/512
  assign sin[337]  =  10'b1100011111;     //337pi/512
  assign cos[337]  =  10'b1110000110;     //337pi/512
  assign sin[338]  =  10'b1100100000;     //338pi/512
  assign cos[338]  =  10'b1110000101;     //338pi/512
  assign sin[339]  =  10'b1100100000;     //339pi/512
  assign cos[339]  =  10'b1110000011;     //339pi/512
  assign sin[340]  =  10'b1100100001;     //340pi/512
  assign cos[340]  =  10'b1110000010;     //340pi/512
  assign sin[341]  =  10'b1100100010;     //341pi/512
  assign cos[341]  =  10'b1110000000;     //341pi/512
  assign sin[342]  =  10'b1100100011;     //342pi/512
  assign cos[342]  =  10'b1101111111;     //342pi/512
  assign sin[343]  =  10'b1100100100;     //343pi/512
  assign cos[343]  =  10'b1101111110;     //343pi/512
  assign sin[344]  =  10'b1100100100;     //344pi/512
  assign cos[344]  =  10'b1101111100;     //344pi/512
  assign sin[345]  =  10'b1100100101;     //345pi/512
  assign cos[345]  =  10'b1101111011;     //345pi/512
  assign sin[346]  =  10'b1100100110;     //346pi/512
  assign cos[346]  =  10'b1101111010;     //346pi/512
  assign sin[347]  =  10'b1100100111;     //347pi/512
  assign cos[347]  =  10'b1101111000;     //347pi/512
  assign sin[348]  =  10'b1100101000;     //348pi/512
  assign cos[348]  =  10'b1101110111;     //348pi/512
  assign sin[349]  =  10'b1100101001;     //349pi/512
  assign cos[349]  =  10'b1101110110;     //349pi/512
  assign sin[350]  =  10'b1100101001;     //350pi/512
  assign cos[350]  =  10'b1101110100;     //350pi/512
  assign sin[351]  =  10'b1100101010;     //351pi/512
  assign cos[351]  =  10'b1101110011;     //351pi/512
  assign sin[352]  =  10'b1100101011;     //352pi/512
  assign cos[352]  =  10'b1101110010;     //352pi/512
  assign sin[353]  =  10'b1100101100;     //353pi/512
  assign cos[353]  =  10'b1101110000;     //353pi/512
  assign sin[354]  =  10'b1100101101;     //354pi/512
  assign cos[354]  =  10'b1101101111;     //354pi/512
  assign sin[355]  =  10'b1100101110;     //355pi/512
  assign cos[355]  =  10'b1101101110;     //355pi/512
  assign sin[356]  =  10'b1100101111;     //356pi/512
  assign cos[356]  =  10'b1101101101;     //356pi/512
  assign sin[357]  =  10'b1100110000;     //357pi/512
  assign cos[357]  =  10'b1101101011;     //357pi/512
  assign sin[358]  =  10'b1100110001;     //358pi/512
  assign cos[358]  =  10'b1101101010;     //358pi/512
  assign sin[359]  =  10'b1100110001;     //359pi/512
  assign cos[359]  =  10'b1101101001;     //359pi/512
  assign sin[360]  =  10'b1100110010;     //360pi/512
  assign cos[360]  =  10'b1101101000;     //360pi/512
  assign sin[361]  =  10'b1100110011;     //361pi/512
  assign cos[361]  =  10'b1101100110;     //361pi/512
  assign sin[362]  =  10'b1100110100;     //362pi/512
  assign cos[362]  =  10'b1101100101;     //362pi/512
  assign sin[363]  =  10'b1100110101;     //363pi/512
  assign cos[363]  =  10'b1101100100;     //363pi/512
  assign sin[364]  =  10'b1100110110;     //364pi/512
  assign cos[364]  =  10'b1101100011;     //364pi/512
  assign sin[365]  =  10'b1100110111;     //365pi/512
  assign cos[365]  =  10'b1101100001;     //365pi/512
  assign sin[366]  =  10'b1100111000;     //366pi/512
  assign cos[366]  =  10'b1101100000;     //366pi/512
  assign sin[367]  =  10'b1100111001;     //367pi/512
  assign cos[367]  =  10'b1101011111;     //367pi/512
  assign sin[368]  =  10'b1100111010;     //368pi/512
  assign cos[368]  =  10'b1101011110;     //368pi/512
  assign sin[369]  =  10'b1100111011;     //369pi/512
  assign cos[369]  =  10'b1101011100;     //369pi/512
  assign sin[370]  =  10'b1100111100;     //370pi/512
  assign cos[370]  =  10'b1101011011;     //370pi/512
  assign sin[371]  =  10'b1100111101;     //371pi/512
  assign cos[371]  =  10'b1101011010;     //371pi/512
  assign sin[372]  =  10'b1100111110;     //372pi/512
  assign cos[372]  =  10'b1101011001;     //372pi/512
  assign sin[373]  =  10'b1100111111;     //373pi/512
  assign cos[373]  =  10'b1101011000;     //373pi/512
  assign sin[374]  =  10'b1101000000;     //374pi/512
  assign cos[374]  =  10'b1101010110;     //374pi/512
  assign sin[375]  =  10'b1101000001;     //375pi/512
  assign cos[375]  =  10'b1101010101;     //375pi/512
  assign sin[376]  =  10'b1101000010;     //376pi/512
  assign cos[376]  =  10'b1101010100;     //376pi/512
  assign sin[377]  =  10'b1101000011;     //377pi/512
  assign cos[377]  =  10'b1101010011;     //377pi/512
  assign sin[378]  =  10'b1101000100;     //378pi/512
  assign cos[378]  =  10'b1101010010;     //378pi/512
  assign sin[379]  =  10'b1101000110;     //379pi/512
  assign cos[379]  =  10'b1101010001;     //379pi/512
  assign sin[380]  =  10'b1101000111;     //380pi/512
  assign cos[380]  =  10'b1101001111;     //380pi/512
  assign sin[381]  =  10'b1101001000;     //381pi/512
  assign cos[381]  =  10'b1101001110;     //381pi/512
  assign sin[382]  =  10'b1101001001;     //382pi/512
  assign cos[382]  =  10'b1101001101;     //382pi/512
  assign sin[383]  =  10'b1101001010;     //383pi/512
  assign cos[383]  =  10'b1101001100;     //383pi/512
  assign sin[384]  =  10'b1101001011;     //384pi/512
  assign cos[384]  =  10'b1101001011;     //384pi/512
  assign sin[385]  =  10'b1101001100;     //385pi/512
  assign cos[385]  =  10'b1101001010;     //385pi/512
  assign sin[386]  =  10'b1101001101;     //386pi/512
  assign cos[386]  =  10'b1101001001;     //386pi/512
  assign sin[387]  =  10'b1101001110;     //387pi/512
  assign cos[387]  =  10'b1101001000;     //387pi/512
  assign sin[388]  =  10'b1101001111;     //388pi/512
  assign cos[388]  =  10'b1101000111;     //388pi/512
  assign sin[389]  =  10'b1101010001;     //389pi/512
  assign cos[389]  =  10'b1101000110;     //389pi/512
  assign sin[390]  =  10'b1101010010;     //390pi/512
  assign cos[390]  =  10'b1101000100;     //390pi/512
  assign sin[391]  =  10'b1101010011;     //391pi/512
  assign cos[391]  =  10'b1101000011;     //391pi/512
  assign sin[392]  =  10'b1101010100;     //392pi/512
  assign cos[392]  =  10'b1101000010;     //392pi/512
  assign sin[393]  =  10'b1101010101;     //393pi/512
  assign cos[393]  =  10'b1101000001;     //393pi/512
  assign sin[394]  =  10'b1101010110;     //394pi/512
  assign cos[394]  =  10'b1101000000;     //394pi/512
  assign sin[395]  =  10'b1101011000;     //395pi/512
  assign cos[395]  =  10'b1100111111;     //395pi/512
  assign sin[396]  =  10'b1101011001;     //396pi/512
  assign cos[396]  =  10'b1100111110;     //396pi/512
  assign sin[397]  =  10'b1101011010;     //397pi/512
  assign cos[397]  =  10'b1100111101;     //397pi/512
  assign sin[398]  =  10'b1101011011;     //398pi/512
  assign cos[398]  =  10'b1100111100;     //398pi/512
  assign sin[399]  =  10'b1101011100;     //399pi/512
  assign cos[399]  =  10'b1100111011;     //399pi/512
  assign sin[400]  =  10'b1101011110;     //400pi/512
  assign cos[400]  =  10'b1100111010;     //400pi/512
  assign sin[401]  =  10'b1101011111;     //401pi/512
  assign cos[401]  =  10'b1100111001;     //401pi/512
  assign sin[402]  =  10'b1101100000;     //402pi/512
  assign cos[402]  =  10'b1100111000;     //402pi/512
  assign sin[403]  =  10'b1101100001;     //403pi/512
  assign cos[403]  =  10'b1100110111;     //403pi/512
  assign sin[404]  =  10'b1101100011;     //404pi/512
  assign cos[404]  =  10'b1100110110;     //404pi/512
  assign sin[405]  =  10'b1101100100;     //405pi/512
  assign cos[405]  =  10'b1100110101;     //405pi/512
  assign sin[406]  =  10'b1101100101;     //406pi/512
  assign cos[406]  =  10'b1100110100;     //406pi/512
  assign sin[407]  =  10'b1101100110;     //407pi/512
  assign cos[407]  =  10'b1100110011;     //407pi/512
  assign sin[408]  =  10'b1101101000;     //408pi/512
  assign cos[408]  =  10'b1100110010;     //408pi/512
  assign sin[409]  =  10'b1101101001;     //409pi/512
  assign cos[409]  =  10'b1100110001;     //409pi/512
  assign sin[410]  =  10'b1101101010;     //410pi/512
  assign cos[410]  =  10'b1100110001;     //410pi/512
  assign sin[411]  =  10'b1101101011;     //411pi/512
  assign cos[411]  =  10'b1100110000;     //411pi/512
  assign sin[412]  =  10'b1101101101;     //412pi/512
  assign cos[412]  =  10'b1100101111;     //412pi/512
  assign sin[413]  =  10'b1101101110;     //413pi/512
  assign cos[413]  =  10'b1100101110;     //413pi/512
  assign sin[414]  =  10'b1101101111;     //414pi/512
  assign cos[414]  =  10'b1100101101;     //414pi/512
  assign sin[415]  =  10'b1101110000;     //415pi/512
  assign cos[415]  =  10'b1100101100;     //415pi/512
  assign sin[416]  =  10'b1101110010;     //416pi/512
  assign cos[416]  =  10'b1100101011;     //416pi/512
  assign sin[417]  =  10'b1101110011;     //417pi/512
  assign cos[417]  =  10'b1100101010;     //417pi/512
  assign sin[418]  =  10'b1101110100;     //418pi/512
  assign cos[418]  =  10'b1100101001;     //418pi/512
  assign sin[419]  =  10'b1101110110;     //419pi/512
  assign cos[419]  =  10'b1100101001;     //419pi/512
  assign sin[420]  =  10'b1101110111;     //420pi/512
  assign cos[420]  =  10'b1100101000;     //420pi/512
  assign sin[421]  =  10'b1101111000;     //421pi/512
  assign cos[421]  =  10'b1100100111;     //421pi/512
  assign sin[422]  =  10'b1101111010;     //422pi/512
  assign cos[422]  =  10'b1100100110;     //422pi/512
  assign sin[423]  =  10'b1101111011;     //423pi/512
  assign cos[423]  =  10'b1100100101;     //423pi/512
  assign sin[424]  =  10'b1101111100;     //424pi/512
  assign cos[424]  =  10'b1100100100;     //424pi/512
  assign sin[425]  =  10'b1101111110;     //425pi/512
  assign cos[425]  =  10'b1100100100;     //425pi/512
  assign sin[426]  =  10'b1101111111;     //426pi/512
  assign cos[426]  =  10'b1100100011;     //426pi/512
  assign sin[427]  =  10'b1110000000;     //427pi/512
  assign cos[427]  =  10'b1100100010;     //427pi/512
  assign sin[428]  =  10'b1110000010;     //428pi/512
  assign cos[428]  =  10'b1100100001;     //428pi/512
  assign sin[429]  =  10'b1110000011;     //429pi/512
  assign cos[429]  =  10'b1100100000;     //429pi/512
  assign sin[430]  =  10'b1110000101;     //430pi/512
  assign cos[430]  =  10'b1100100000;     //430pi/512
  assign sin[431]  =  10'b1110000110;     //431pi/512
  assign cos[431]  =  10'b1100011111;     //431pi/512
  assign sin[432]  =  10'b1110000111;     //432pi/512
  assign cos[432]  =  10'b1100011110;     //432pi/512
  assign sin[433]  =  10'b1110001001;     //433pi/512
  assign cos[433]  =  10'b1100011101;     //433pi/512
  assign sin[434]  =  10'b1110001010;     //434pi/512
  assign cos[434]  =  10'b1100011101;     //434pi/512
  assign sin[435]  =  10'b1110001011;     //435pi/512
  assign cos[435]  =  10'b1100011100;     //435pi/512
  assign sin[436]  =  10'b1110001101;     //436pi/512
  assign cos[436]  =  10'b1100011011;     //436pi/512
  assign sin[437]  =  10'b1110001110;     //437pi/512
  assign cos[437]  =  10'b1100011011;     //437pi/512
  assign sin[438]  =  10'b1110010000;     //438pi/512
  assign cos[438]  =  10'b1100011010;     //438pi/512
  assign sin[439]  =  10'b1110010001;     //439pi/512
  assign cos[439]  =  10'b1100011001;     //439pi/512
  assign sin[440]  =  10'b1110010011;     //440pi/512
  assign cos[440]  =  10'b1100011001;     //440pi/512
  assign sin[441]  =  10'b1110010100;     //441pi/512
  assign cos[441]  =  10'b1100011000;     //441pi/512
  assign sin[442]  =  10'b1110010101;     //442pi/512
  assign cos[442]  =  10'b1100010111;     //442pi/512
  assign sin[443]  =  10'b1110010111;     //443pi/512
  assign cos[443]  =  10'b1100010111;     //443pi/512
  assign sin[444]  =  10'b1110011000;     //444pi/512
  assign cos[444]  =  10'b1100010110;     //444pi/512
  assign sin[445]  =  10'b1110011010;     //445pi/512
  assign cos[445]  =  10'b1100010101;     //445pi/512
  assign sin[446]  =  10'b1110011011;     //446pi/512
  assign cos[446]  =  10'b1100010101;     //446pi/512
  assign sin[447]  =  10'b1110011101;     //447pi/512
  assign cos[447]  =  10'b1100010100;     //447pi/512
  assign sin[448]  =  10'b1110011110;     //448pi/512
  assign cos[448]  =  10'b1100010011;     //448pi/512
  assign sin[449]  =  10'b1110011111;     //449pi/512
  assign cos[449]  =  10'b1100010011;     //449pi/512
  assign sin[450]  =  10'b1110100001;     //450pi/512
  assign cos[450]  =  10'b1100010010;     //450pi/512
  assign sin[451]  =  10'b1110100010;     //451pi/512
  assign cos[451]  =  10'b1100010010;     //451pi/512
  assign sin[452]  =  10'b1110100100;     //452pi/512
  assign cos[452]  =  10'b1100010001;     //452pi/512
  assign sin[453]  =  10'b1110100101;     //453pi/512
  assign cos[453]  =  10'b1100010001;     //453pi/512
  assign sin[454]  =  10'b1110100111;     //454pi/512
  assign cos[454]  =  10'b1100010000;     //454pi/512
  assign sin[455]  =  10'b1110101000;     //455pi/512
  assign cos[455]  =  10'b1100001111;     //455pi/512
  assign sin[456]  =  10'b1110101010;     //456pi/512
  assign cos[456]  =  10'b1100001111;     //456pi/512
  assign sin[457]  =  10'b1110101011;     //457pi/512
  assign cos[457]  =  10'b1100001110;     //457pi/512
  assign sin[458]  =  10'b1110101101;     //458pi/512
  assign cos[458]  =  10'b1100001110;     //458pi/512
  assign sin[459]  =  10'b1110101110;     //459pi/512
  assign cos[459]  =  10'b1100001101;     //459pi/512
  assign sin[460]  =  10'b1110110000;     //460pi/512
  assign cos[460]  =  10'b1100001101;     //460pi/512
  assign sin[461]  =  10'b1110110001;     //461pi/512
  assign cos[461]  =  10'b1100001100;     //461pi/512
  assign sin[462]  =  10'b1110110011;     //462pi/512
  assign cos[462]  =  10'b1100001100;     //462pi/512
  assign sin[463]  =  10'b1110110100;     //463pi/512
  assign cos[463]  =  10'b1100001011;     //463pi/512
  assign sin[464]  =  10'b1110110110;     //464pi/512
  assign cos[464]  =  10'b1100001011;     //464pi/512
  assign sin[465]  =  10'b1110110111;     //465pi/512
  assign cos[465]  =  10'b1100001011;     //465pi/512
  assign sin[466]  =  10'b1110111001;     //466pi/512
  assign cos[466]  =  10'b1100001010;     //466pi/512
  assign sin[467]  =  10'b1110111010;     //467pi/512
  assign cos[467]  =  10'b1100001010;     //467pi/512
  assign sin[468]  =  10'b1110111100;     //468pi/512
  assign cos[468]  =  10'b1100001001;     //468pi/512
  assign sin[469]  =  10'b1110111101;     //469pi/512
  assign cos[469]  =  10'b1100001001;     //469pi/512
  assign sin[470]  =  10'b1110111111;     //470pi/512
  assign cos[470]  =  10'b1100001000;     //470pi/512
  assign sin[471]  =  10'b1111000000;     //471pi/512
  assign cos[471]  =  10'b1100001000;     //471pi/512
  assign sin[472]  =  10'b1111000010;     //472pi/512
  assign cos[472]  =  10'b1100001000;     //472pi/512
  assign sin[473]  =  10'b1111000011;     //473pi/512
  assign cos[473]  =  10'b1100000111;     //473pi/512
  assign sin[474]  =  10'b1111000101;     //474pi/512
  assign cos[474]  =  10'b1100000111;     //474pi/512
  assign sin[475]  =  10'b1111000110;     //475pi/512
  assign cos[475]  =  10'b1100000111;     //475pi/512
  assign sin[476]  =  10'b1111001000;     //476pi/512
  assign cos[476]  =  10'b1100000110;     //476pi/512
  assign sin[477]  =  10'b1111001001;     //477pi/512
  assign cos[477]  =  10'b1100000110;     //477pi/512
  assign sin[478]  =  10'b1111001011;     //478pi/512
  assign cos[478]  =  10'b1100000110;     //478pi/512
  assign sin[479]  =  10'b1111001101;     //479pi/512
  assign cos[479]  =  10'b1100000101;     //479pi/512
  assign sin[480]  =  10'b1111001110;     //480pi/512
  assign cos[480]  =  10'b1100000101;     //480pi/512
  assign sin[481]  =  10'b1111010000;     //481pi/512
  assign cos[481]  =  10'b1100000101;     //481pi/512
  assign sin[482]  =  10'b1111010001;     //482pi/512
  assign cos[482]  =  10'b1100000100;     //482pi/512
  assign sin[483]  =  10'b1111010011;     //483pi/512
  assign cos[483]  =  10'b1100000100;     //483pi/512
  assign sin[484]  =  10'b1111010100;     //484pi/512
  assign cos[484]  =  10'b1100000100;     //484pi/512
  assign sin[485]  =  10'b1111010110;     //485pi/512
  assign cos[485]  =  10'b1100000100;     //485pi/512
  assign sin[486]  =  10'b1111010111;     //486pi/512
  assign cos[486]  =  10'b1100000011;     //486pi/512
  assign sin[487]  =  10'b1111011001;     //487pi/512
  assign cos[487]  =  10'b1100000011;     //487pi/512
  assign sin[488]  =  10'b1111011010;     //488pi/512
  assign cos[488]  =  10'b1100000011;     //488pi/512
  assign sin[489]  =  10'b1111011100;     //489pi/512
  assign cos[489]  =  10'b1100000011;     //489pi/512
  assign sin[490]  =  10'b1111011110;     //490pi/512
  assign cos[490]  =  10'b1100000010;     //490pi/512
  assign sin[491]  =  10'b1111011111;     //491pi/512
  assign cos[491]  =  10'b1100000010;     //491pi/512
  assign sin[492]  =  10'b1111100001;     //492pi/512
  assign cos[492]  =  10'b1100000010;     //492pi/512
  assign sin[493]  =  10'b1111100010;     //493pi/512
  assign cos[493]  =  10'b1100000010;     //493pi/512
  assign sin[494]  =  10'b1111100100;     //494pi/512
  assign cos[494]  =  10'b1100000010;     //494pi/512
  assign sin[495]  =  10'b1111100101;     //495pi/512
  assign cos[495]  =  10'b1100000001;     //495pi/512
  assign sin[496]  =  10'b1111100111;     //496pi/512
  assign cos[496]  =  10'b1100000001;     //496pi/512
  assign sin[497]  =  10'b1111101000;     //497pi/512
  assign cos[497]  =  10'b1100000001;     //497pi/512
  assign sin[498]  =  10'b1111101010;     //498pi/512
  assign cos[498]  =  10'b1100000001;     //498pi/512
  assign sin[499]  =  10'b1111101100;     //499pi/512
  assign cos[499]  =  10'b1100000001;     //499pi/512
  assign sin[500]  =  10'b1111101101;     //500pi/512
  assign cos[500]  =  10'b1100000001;     //500pi/512
  assign sin[501]  =  10'b1111101111;     //501pi/512
  assign cos[501]  =  10'b1100000001;     //501pi/512
  assign sin[502]  =  10'b1111110000;     //502pi/512
  assign cos[502]  =  10'b1100000000;     //502pi/512
  assign sin[503]  =  10'b1111110010;     //503pi/512
  assign cos[503]  =  10'b1100000000;     //503pi/512
  assign sin[504]  =  10'b1111110011;     //504pi/512
  assign cos[504]  =  10'b1100000000;     //504pi/512
  assign sin[505]  =  10'b1111110101;     //505pi/512
  assign cos[505]  =  10'b1100000000;     //505pi/512
  assign sin[506]  =  10'b1111110111;     //506pi/512
  assign cos[506]  =  10'b1100000000;     //506pi/512
  assign sin[507]  =  10'b1111111000;     //507pi/512
  assign cos[507]  =  10'b1100000000;     //507pi/512
  assign sin[508]  =  10'b1111111010;     //508pi/512
  assign cos[508]  =  10'b1100000000;     //508pi/512
  assign sin[509]  =  10'b1111111011;     //509pi/512
  assign cos[509]  =  10'b1100000000;     //509pi/512
  assign sin[510]  =  10'b1111111101;     //510pi/512
  assign cos[510]  =  10'b1100000000;     //510pi/512
  assign sin[511]  =  10'b1111111110;     //511pi/512
  assign cos[511]  =  10'b1100000000;     //511pi/512
endmodule