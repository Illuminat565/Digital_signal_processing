module  TWIDLE_14_bit  #(parameter stage_FFT = 2, SIZE =10, word_length_tw = 14) (
    input            clk,
    input            en_rd, 
    input   [stage_FFT-2:0]   rd_ptr_angle,

    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );

reg signed [word_length_tw-1:0]  cos  [511:0];
reg signed [word_length_tw-1:0]  sin  [511:0];

//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd) begin
                  cos_data           <= cos   [rd_ptr_angle];
                  sin_data           <= sin   [rd_ptr_angle];
             end 
        end
//----------------------------------------------------------------------------------------
initial begin
   sin[0]  =  14'b00000000000000;     //0pi/1024
   cos[0]  =  14'b01000000000000;     //0pi/1024
   sin[1]  =  14'b11111111100111;     //2pi/1024
   cos[1]  =  14'b00111111111111;     //2pi/1024
   sin[2]  =  14'b11111111001110;     //4pi/1024
   cos[2]  =  14'b00111111111111;     //4pi/1024
   sin[3]  =  14'b11111110110101;     //6pi/1024
   cos[3]  =  14'b00111111111111;     //6pi/1024
   sin[4]  =  14'b11111110011011;     //8pi/1024
   cos[4]  =  14'b00111111111110;     //8pi/1024
   sin[5]  =  14'b11111110000010;     //10pi/1024
   cos[5]  =  14'b00111111111110;     //10pi/1024
   sin[6]  =  14'b11111101101001;     //12pi/1024
   cos[6]  =  14'b00111111111101;     //12pi/1024
   sin[7]  =  14'b11111101010000;     //14pi/1024
   cos[7]  =  14'b00111111111100;     //14pi/1024
   sin[8]  =  14'b11111100110111;     //16pi/1024
   cos[8]  =  14'b00111111111011;     //16pi/1024
   sin[9]  =  14'b11111100011110;     //18pi/1024
   cos[9]  =  14'b00111111111001;     //18pi/1024
   sin[10]  =  14'b11111100000101;     //20pi/1024
   cos[10]  =  14'b00111111111000;     //20pi/1024
   sin[11]  =  14'b11111011101100;     //22pi/1024
   cos[11]  =  14'b00111111110110;     //22pi/1024
   sin[12]  =  14'b11111011010011;     //24pi/1024
   cos[12]  =  14'b00111111110100;     //24pi/1024
   sin[13]  =  14'b11111010111010;     //26pi/1024
   cos[13]  =  14'b00111111110010;     //26pi/1024
   sin[14]  =  14'b11111010100001;     //28pi/1024
   cos[14]  =  14'b00111111110000;     //28pi/1024
   sin[15]  =  14'b11111010001000;     //30pi/1024
   cos[15]  =  14'b00111111101110;     //30pi/1024
   sin[16]  =  14'b11111001101111;     //32pi/1024
   cos[16]  =  14'b00111111101100;     //32pi/1024
   sin[17]  =  14'b11111001010110;     //34pi/1024
   cos[17]  =  14'b00111111101001;     //34pi/1024
   sin[18]  =  14'b11111000111101;     //36pi/1024
   cos[18]  =  14'b00111111100111;     //36pi/1024
   sin[19]  =  14'b11111000100100;     //38pi/1024
   cos[19]  =  14'b00111111100100;     //38pi/1024
   sin[20]  =  14'b11111000001011;     //40pi/1024
   cos[20]  =  14'b00111111100001;     //40pi/1024
   sin[21]  =  14'b11110111110010;     //42pi/1024
   cos[21]  =  14'b00111111011110;     //42pi/1024
   sin[22]  =  14'b11110111011001;     //44pi/1024
   cos[22]  =  14'b00111111011010;     //44pi/1024
   sin[23]  =  14'b11110111000000;     //46pi/1024
   cos[23]  =  14'b00111111010111;     //46pi/1024
   sin[24]  =  14'b11110110100111;     //48pi/1024
   cos[24]  =  14'b00111111010011;     //48pi/1024
   sin[25]  =  14'b11110110001110;     //50pi/1024
   cos[25]  =  14'b00111111001111;     //50pi/1024
   sin[26]  =  14'b11110101110101;     //52pi/1024
   cos[26]  =  14'b00111111001011;     //52pi/1024
   sin[27]  =  14'b11110101011101;     //54pi/1024
   cos[27]  =  14'b00111111000111;     //54pi/1024
   sin[28]  =  14'b11110101000100;     //56pi/1024
   cos[28]  =  14'b00111111000011;     //56pi/1024
   sin[29]  =  14'b11110100101011;     //58pi/1024
   cos[29]  =  14'b00111110111111;     //58pi/1024
   sin[30]  =  14'b11110100010010;     //60pi/1024
   cos[30]  =  14'b00111110111010;     //60pi/1024
   sin[31]  =  14'b11110011111010;     //62pi/1024
   cos[31]  =  14'b00111110110110;     //62pi/1024
   sin[32]  =  14'b11110011100001;     //64pi/1024
   cos[32]  =  14'b00111110110001;     //64pi/1024
   sin[33]  =  14'b11110011001000;     //66pi/1024
   cos[33]  =  14'b00111110101100;     //66pi/1024
   sin[34]  =  14'b11110010110000;     //68pi/1024
   cos[34]  =  14'b00111110100111;     //68pi/1024
   sin[35]  =  14'b11110010010111;     //70pi/1024
   cos[35]  =  14'b00111110100001;     //70pi/1024
   sin[36]  =  14'b11110001111111;     //72pi/1024
   cos[36]  =  14'b00111110011100;     //72pi/1024
   sin[37]  =  14'b11110001100110;     //74pi/1024
   cos[37]  =  14'b00111110010110;     //74pi/1024
   sin[38]  =  14'b11110001001110;     //76pi/1024
   cos[38]  =  14'b00111110010001;     //76pi/1024
   sin[39]  =  14'b11110000110101;     //78pi/1024
   cos[39]  =  14'b00111110001011;     //78pi/1024
   sin[40]  =  14'b11110000011101;     //80pi/1024
   cos[40]  =  14'b00111110000101;     //80pi/1024
   sin[41]  =  14'b11110000000100;     //82pi/1024
   cos[41]  =  14'b00111101111111;     //82pi/1024
   sin[42]  =  14'b11101111101100;     //84pi/1024
   cos[42]  =  14'b00111101111000;     //84pi/1024
   sin[43]  =  14'b11101111010100;     //86pi/1024
   cos[43]  =  14'b00111101110010;     //86pi/1024
   sin[44]  =  14'b11101110111100;     //88pi/1024
   cos[44]  =  14'b00111101101011;     //88pi/1024
   sin[45]  =  14'b11101110100011;     //90pi/1024
   cos[45]  =  14'b00111101100100;     //90pi/1024
   sin[46]  =  14'b11101110001011;     //92pi/1024
   cos[46]  =  14'b00111101011101;     //92pi/1024
   sin[47]  =  14'b11101101110011;     //94pi/1024
   cos[47]  =  14'b00111101010110;     //94pi/1024
   sin[48]  =  14'b11101101011011;     //96pi/1024
   cos[48]  =  14'b00111101001111;     //96pi/1024
   sin[49]  =  14'b11101101000011;     //98pi/1024
   cos[49]  =  14'b00111101001000;     //98pi/1024
   sin[50]  =  14'b11101100101011;     //100pi/1024
   cos[50]  =  14'b00111101000000;     //100pi/1024
   sin[51]  =  14'b11101100010011;     //102pi/1024
   cos[51]  =  14'b00111100111001;     //102pi/1024
   sin[52]  =  14'b11101011111011;     //104pi/1024
   cos[52]  =  14'b00111100110001;     //104pi/1024
   sin[53]  =  14'b11101011100011;     //106pi/1024
   cos[53]  =  14'b00111100101001;     //106pi/1024
   sin[54]  =  14'b11101011001100;     //108pi/1024
   cos[54]  =  14'b00111100100001;     //108pi/1024
   sin[55]  =  14'b11101010110100;     //110pi/1024
   cos[55]  =  14'b00111100011000;     //110pi/1024
   sin[56]  =  14'b11101010011100;     //112pi/1024
   cos[56]  =  14'b00111100010000;     //112pi/1024
   sin[57]  =  14'b11101010000100;     //114pi/1024
   cos[57]  =  14'b00111100001000;     //114pi/1024
   sin[58]  =  14'b11101001101101;     //116pi/1024
   cos[58]  =  14'b00111011111111;     //116pi/1024
   sin[59]  =  14'b11101001010101;     //118pi/1024
   cos[59]  =  14'b00111011110110;     //118pi/1024
   sin[60]  =  14'b11101000111110;     //120pi/1024
   cos[60]  =  14'b00111011101101;     //120pi/1024
   sin[61]  =  14'b11101000100110;     //122pi/1024
   cos[61]  =  14'b00111011100100;     //122pi/1024
   sin[62]  =  14'b11101000001111;     //124pi/1024
   cos[62]  =  14'b00111011011011;     //124pi/1024
   sin[63]  =  14'b11100111111000;     //126pi/1024
   cos[63]  =  14'b00111011010001;     //126pi/1024
   sin[64]  =  14'b11100111100001;     //128pi/1024
   cos[64]  =  14'b00111011001000;     //128pi/1024
   sin[65]  =  14'b11100111001001;     //130pi/1024
   cos[65]  =  14'b00111010111110;     //130pi/1024
   sin[66]  =  14'b11100110110010;     //132pi/1024
   cos[66]  =  14'b00111010110100;     //132pi/1024
   sin[67]  =  14'b11100110011011;     //134pi/1024
   cos[67]  =  14'b00111010101010;     //134pi/1024
   sin[68]  =  14'b11100110000100;     //136pi/1024
   cos[68]  =  14'b00111010100000;     //136pi/1024
   sin[69]  =  14'b11100101101101;     //138pi/1024
   cos[69]  =  14'b00111010010110;     //138pi/1024
   sin[70]  =  14'b11100101010110;     //140pi/1024
   cos[70]  =  14'b00111010001011;     //140pi/1024
   sin[71]  =  14'b11100100111111;     //142pi/1024
   cos[71]  =  14'b00111010000001;     //142pi/1024
   sin[72]  =  14'b11100100101001;     //144pi/1024
   cos[72]  =  14'b00111001110110;     //144pi/1024
   sin[73]  =  14'b11100100010010;     //146pi/1024
   cos[73]  =  14'b00111001101011;     //146pi/1024
   sin[74]  =  14'b11100011111011;     //148pi/1024
   cos[74]  =  14'b00111001100000;     //148pi/1024
   sin[75]  =  14'b11100011100101;     //150pi/1024
   cos[75]  =  14'b00111001010101;     //150pi/1024
   sin[76]  =  14'b11100011001110;     //152pi/1024
   cos[76]  =  14'b00111001001010;     //152pi/1024
   sin[77]  =  14'b11100010111000;     //154pi/1024
   cos[77]  =  14'b00111000111111;     //154pi/1024
   sin[78]  =  14'b11100010100010;     //156pi/1024
   cos[78]  =  14'b00111000110011;     //156pi/1024
   sin[79]  =  14'b11100010001011;     //158pi/1024
   cos[79]  =  14'b00111000101000;     //158pi/1024
   sin[80]  =  14'b11100001110101;     //160pi/1024
   cos[80]  =  14'b00111000011100;     //160pi/1024
   sin[81]  =  14'b11100001011111;     //162pi/1024
   cos[81]  =  14'b00111000010000;     //162pi/1024
   sin[82]  =  14'b11100001001001;     //164pi/1024
   cos[82]  =  14'b00111000000100;     //164pi/1024
   sin[83]  =  14'b11100000110011;     //166pi/1024
   cos[83]  =  14'b00110111111000;     //166pi/1024
   sin[84]  =  14'b11100000011101;     //168pi/1024
   cos[84]  =  14'b00110111101011;     //168pi/1024
   sin[85]  =  14'b11100000000111;     //170pi/1024
   cos[85]  =  14'b00110111011111;     //170pi/1024
   sin[86]  =  14'b11011111110010;     //172pi/1024
   cos[86]  =  14'b00110111010010;     //172pi/1024
   sin[87]  =  14'b11011111011100;     //174pi/1024
   cos[87]  =  14'b00110111000110;     //174pi/1024
   sin[88]  =  14'b11011111000110;     //176pi/1024
   cos[88]  =  14'b00110110111001;     //176pi/1024
   sin[89]  =  14'b11011110110001;     //178pi/1024
   cos[89]  =  14'b00110110101100;     //178pi/1024
   sin[90]  =  14'b11011110011011;     //180pi/1024
   cos[90]  =  14'b00110110011111;     //180pi/1024
   sin[91]  =  14'b11011110000110;     //182pi/1024
   cos[91]  =  14'b00110110010001;     //182pi/1024
   sin[92]  =  14'b11011101110001;     //184pi/1024
   cos[92]  =  14'b00110110000100;     //184pi/1024
   sin[93]  =  14'b11011101011011;     //186pi/1024
   cos[93]  =  14'b00110101110111;     //186pi/1024
   sin[94]  =  14'b11011101000110;     //188pi/1024
   cos[94]  =  14'b00110101101001;     //188pi/1024
   sin[95]  =  14'b11011100110001;     //190pi/1024
   cos[95]  =  14'b00110101011011;     //190pi/1024
   sin[96]  =  14'b11011100011100;     //192pi/1024
   cos[96]  =  14'b00110101001101;     //192pi/1024
   sin[97]  =  14'b11011100001000;     //194pi/1024
   cos[97]  =  14'b00110100111111;     //194pi/1024
   sin[98]  =  14'b11011011110011;     //196pi/1024
   cos[98]  =  14'b00110100110001;     //196pi/1024
   sin[99]  =  14'b11011011011110;     //198pi/1024
   cos[99]  =  14'b00110100100011;     //198pi/1024
   sin[100]  =  14'b11011011001001;     //200pi/1024
   cos[100]  =  14'b00110100010100;     //200pi/1024
   sin[101]  =  14'b11011010110101;     //202pi/1024
   cos[101]  =  14'b00110100000110;     //202pi/1024
   sin[102]  =  14'b11011010100001;     //204pi/1024
   cos[102]  =  14'b00110011110111;     //204pi/1024
   sin[103]  =  14'b11011010001100;     //206pi/1024
   cos[103]  =  14'b00110011101000;     //206pi/1024
   sin[104]  =  14'b11011001111000;     //208pi/1024
   cos[104]  =  14'b00110011011001;     //208pi/1024
   sin[105]  =  14'b11011001100100;     //210pi/1024
   cos[105]  =  14'b00110011001010;     //210pi/1024
   sin[106]  =  14'b11011001010000;     //212pi/1024
   cos[106]  =  14'b00110010111011;     //212pi/1024
   sin[107]  =  14'b11011000111100;     //214pi/1024
   cos[107]  =  14'b00110010101100;     //214pi/1024
   sin[108]  =  14'b11011000101000;     //216pi/1024
   cos[108]  =  14'b00110010011101;     //216pi/1024
   sin[109]  =  14'b11011000010100;     //218pi/1024
   cos[109]  =  14'b00110010001101;     //218pi/1024
   sin[110]  =  14'b11011000000001;     //220pi/1024
   cos[110]  =  14'b00110001111101;     //220pi/1024
   sin[111]  =  14'b11010111101101;     //222pi/1024
   cos[111]  =  14'b00110001101110;     //222pi/1024
   sin[112]  =  14'b11010111011010;     //224pi/1024
   cos[112]  =  14'b00110001011110;     //224pi/1024
   sin[113]  =  14'b11010111000110;     //226pi/1024
   cos[113]  =  14'b00110001001110;     //226pi/1024
   sin[114]  =  14'b11010110110011;     //228pi/1024
   cos[114]  =  14'b00110000111110;     //228pi/1024
   sin[115]  =  14'b11010110100000;     //230pi/1024
   cos[115]  =  14'b00110000101101;     //230pi/1024
   sin[116]  =  14'b11010110001101;     //232pi/1024
   cos[116]  =  14'b00110000011101;     //232pi/1024
   sin[117]  =  14'b11010101111010;     //234pi/1024
   cos[117]  =  14'b00110000001101;     //234pi/1024
   sin[118]  =  14'b11010101100111;     //236pi/1024
   cos[118]  =  14'b00101111111100;     //236pi/1024
   sin[119]  =  14'b11010101010100;     //238pi/1024
   cos[119]  =  14'b00101111101011;     //238pi/1024
   sin[120]  =  14'b11010101000001;     //240pi/1024
   cos[120]  =  14'b00101111011010;     //240pi/1024
   sin[121]  =  14'b11010100101111;     //242pi/1024
   cos[121]  =  14'b00101111001010;     //242pi/1024
   sin[122]  =  14'b11010100011100;     //244pi/1024
   cos[122]  =  14'b00101110111000;     //244pi/1024
   sin[123]  =  14'b11010100001010;     //246pi/1024
   cos[123]  =  14'b00101110100111;     //246pi/1024
   sin[124]  =  14'b11010011111000;     //248pi/1024
   cos[124]  =  14'b00101110010110;     //248pi/1024
   sin[125]  =  14'b11010011100101;     //250pi/1024
   cos[125]  =  14'b00101110000101;     //250pi/1024
   sin[126]  =  14'b11010011010011;     //252pi/1024
   cos[126]  =  14'b00101101110011;     //252pi/1024
   sin[127]  =  14'b11010011000010;     //254pi/1024
   cos[127]  =  14'b00101101100010;     //254pi/1024
   sin[128]  =  14'b11010010110000;     //256pi/1024
   cos[128]  =  14'b00101101010000;     //256pi/1024
   sin[129]  =  14'b11010010011110;     //258pi/1024
   cos[129]  =  14'b00101100111110;     //258pi/1024
   sin[130]  =  14'b11010010001100;     //260pi/1024
   cos[130]  =  14'b00101100101100;     //260pi/1024
   sin[131]  =  14'b11010001111011;     //262pi/1024
   cos[131]  =  14'b00101100011010;     //262pi/1024
   sin[132]  =  14'b11010001101001;     //264pi/1024
   cos[132]  =  14'b00101100001000;     //264pi/1024
   sin[133]  =  14'b11010001011000;     //266pi/1024
   cos[133]  =  14'b00101011110110;     //266pi/1024
   sin[134]  =  14'b11010001000111;     //268pi/1024
   cos[134]  =  14'b00101011100011;     //268pi/1024
   sin[135]  =  14'b11010000110110;     //270pi/1024
   cos[135]  =  14'b00101011010001;     //270pi/1024
   sin[136]  =  14'b11010000100101;     //272pi/1024
   cos[136]  =  14'b00101010111110;     //272pi/1024
   sin[137]  =  14'b11010000010100;     //274pi/1024
   cos[137]  =  14'b00101010101100;     //274pi/1024
   sin[138]  =  14'b11010000000100;     //276pi/1024
   cos[138]  =  14'b00101010011001;     //276pi/1024
   sin[139]  =  14'b11001111110011;     //278pi/1024
   cos[139]  =  14'b00101010000110;     //278pi/1024
   sin[140]  =  14'b11001111100010;     //280pi/1024
   cos[140]  =  14'b00101001110011;     //280pi/1024
   sin[141]  =  14'b11001111010010;     //282pi/1024
   cos[141]  =  14'b00101001100000;     //282pi/1024
   sin[142]  =  14'b11001111000010;     //284pi/1024
   cos[142]  =  14'b00101001001101;     //284pi/1024
   sin[143]  =  14'b11001110110010;     //286pi/1024
   cos[143]  =  14'b00101000111001;     //286pi/1024
   sin[144]  =  14'b11001110100010;     //288pi/1024
   cos[144]  =  14'b00101000100110;     //288pi/1024
   sin[145]  =  14'b11001110010010;     //290pi/1024
   cos[145]  =  14'b00101000010010;     //290pi/1024
   sin[146]  =  14'b11001110000010;     //292pi/1024
   cos[146]  =  14'b00100111111111;     //292pi/1024
   sin[147]  =  14'b11001101110010;     //294pi/1024
   cos[147]  =  14'b00100111101011;     //294pi/1024
   sin[148]  =  14'b11001101100011;     //296pi/1024
   cos[148]  =  14'b00100111010111;     //296pi/1024
   sin[149]  =  14'b11001101010100;     //298pi/1024
   cos[149]  =  14'b00100111000100;     //298pi/1024
   sin[150]  =  14'b11001101000100;     //300pi/1024
   cos[150]  =  14'b00100110110000;     //300pi/1024
   sin[151]  =  14'b11001100110101;     //302pi/1024
   cos[151]  =  14'b00100110011100;     //302pi/1024
   sin[152]  =  14'b11001100100110;     //304pi/1024
   cos[152]  =  14'b00100110000111;     //304pi/1024
   sin[153]  =  14'b11001100010111;     //306pi/1024
   cos[153]  =  14'b00100101110011;     //306pi/1024
   sin[154]  =  14'b11001100001000;     //308pi/1024
   cos[154]  =  14'b00100101011111;     //308pi/1024
   sin[155]  =  14'b11001011111010;     //310pi/1024
   cos[155]  =  14'b00100101001011;     //310pi/1024
   sin[156]  =  14'b11001011101011;     //312pi/1024
   cos[156]  =  14'b00100100110110;     //312pi/1024
   sin[157]  =  14'b11001011011101;     //314pi/1024
   cos[157]  =  14'b00100100100001;     //314pi/1024
   sin[158]  =  14'b11001011001110;     //316pi/1024
   cos[158]  =  14'b00100100001101;     //316pi/1024
   sin[159]  =  14'b11001011000000;     //318pi/1024
   cos[159]  =  14'b00100011111000;     //318pi/1024
   sin[160]  =  14'b11001010110010;     //320pi/1024
   cos[160]  =  14'b00100011100011;     //320pi/1024
   sin[161]  =  14'b11001010100100;     //322pi/1024
   cos[161]  =  14'b00100011001110;     //322pi/1024
   sin[162]  =  14'b11001010010111;     //324pi/1024
   cos[162]  =  14'b00100010111001;     //324pi/1024
   sin[163]  =  14'b11001010001001;     //326pi/1024
   cos[163]  =  14'b00100010100100;     //326pi/1024
   sin[164]  =  14'b11001001111011;     //328pi/1024
   cos[164]  =  14'b00100010001111;     //328pi/1024
   sin[165]  =  14'b11001001101110;     //330pi/1024
   cos[165]  =  14'b00100001111010;     //330pi/1024
   sin[166]  =  14'b11001001100001;     //332pi/1024
   cos[166]  =  14'b00100001100100;     //332pi/1024
   sin[167]  =  14'b11001001010100;     //334pi/1024
   cos[167]  =  14'b00100001001111;     //334pi/1024
   sin[168]  =  14'b11001001000111;     //336pi/1024
   cos[168]  =  14'b00100000111001;     //336pi/1024
   sin[169]  =  14'b11001000111010;     //338pi/1024
   cos[169]  =  14'b00100000100100;     //338pi/1024
   sin[170]  =  14'b11001000101101;     //340pi/1024
   cos[170]  =  14'b00100000001110;     //340pi/1024
   sin[171]  =  14'b11001000100001;     //342pi/1024
   cos[171]  =  14'b00011111111000;     //342pi/1024
   sin[172]  =  14'b11001000010100;     //344pi/1024
   cos[172]  =  14'b00011111100010;     //344pi/1024
   sin[173]  =  14'b11001000001000;     //346pi/1024
   cos[173]  =  14'b00011111001101;     //346pi/1024
   sin[174]  =  14'b11000111111100;     //348pi/1024
   cos[174]  =  14'b00011110110111;     //348pi/1024
   sin[175]  =  14'b11000111110000;     //350pi/1024
   cos[175]  =  14'b00011110100000;     //350pi/1024
   sin[176]  =  14'b11000111100100;     //352pi/1024
   cos[176]  =  14'b00011110001010;     //352pi/1024
   sin[177]  =  14'b11000111011000;     //354pi/1024
   cos[177]  =  14'b00011101110100;     //354pi/1024
   sin[178]  =  14'b11000111001100;     //356pi/1024
   cos[178]  =  14'b00011101011110;     //356pi/1024
   sin[179]  =  14'b11000111000001;     //358pi/1024
   cos[179]  =  14'b00011101001000;     //358pi/1024
   sin[180]  =  14'b11000110110101;     //360pi/1024
   cos[180]  =  14'b00011100110001;     //360pi/1024
   sin[181]  =  14'b11000110101010;     //362pi/1024
   cos[181]  =  14'b00011100011011;     //362pi/1024
   sin[182]  =  14'b11000110011111;     //364pi/1024
   cos[182]  =  14'b00011100000100;     //364pi/1024
   sin[183]  =  14'b11000110010100;     //366pi/1024
   cos[183]  =  14'b00011011101101;     //366pi/1024
   sin[184]  =  14'b11000110001001;     //368pi/1024
   cos[184]  =  14'b00011011010111;     //368pi/1024
   sin[185]  =  14'b11000101111111;     //370pi/1024
   cos[185]  =  14'b00011011000000;     //370pi/1024
   sin[186]  =  14'b11000101110100;     //372pi/1024
   cos[186]  =  14'b00011010101001;     //372pi/1024
   sin[187]  =  14'b11000101101010;     //374pi/1024
   cos[187]  =  14'b00011010010010;     //374pi/1024
   sin[188]  =  14'b11000101011111;     //376pi/1024
   cos[188]  =  14'b00011001111011;     //376pi/1024
   sin[189]  =  14'b11000101010101;     //378pi/1024
   cos[189]  =  14'b00011001100100;     //378pi/1024
   sin[190]  =  14'b11000101001011;     //380pi/1024
   cos[190]  =  14'b00011001001101;     //380pi/1024
   sin[191]  =  14'b11000101000001;     //382pi/1024
   cos[191]  =  14'b00011000110110;     //382pi/1024
   sin[192]  =  14'b11000100111000;     //384pi/1024
   cos[192]  =  14'b00011000011111;     //384pi/1024
   sin[193]  =  14'b11000100101110;     //386pi/1024
   cos[193]  =  14'b00011000001000;     //386pi/1024
   sin[194]  =  14'b11000100100101;     //388pi/1024
   cos[194]  =  14'b00010111110000;     //388pi/1024
   sin[195]  =  14'b11000100011100;     //390pi/1024
   cos[195]  =  14'b00010111011001;     //390pi/1024
   sin[196]  =  14'b11000100010010;     //392pi/1024
   cos[196]  =  14'b00010111000010;     //392pi/1024
   sin[197]  =  14'b11000100001001;     //394pi/1024
   cos[197]  =  14'b00010110101010;     //394pi/1024
   sin[198]  =  14'b11000100000001;     //396pi/1024
   cos[198]  =  14'b00010110010011;     //396pi/1024
   sin[199]  =  14'b11000011111000;     //398pi/1024
   cos[199]  =  14'b00010101111011;     //398pi/1024
   sin[200]  =  14'b11000011101111;     //400pi/1024
   cos[200]  =  14'b00010101100011;     //400pi/1024
   sin[201]  =  14'b11000011100111;     //402pi/1024
   cos[201]  =  14'b00010101001100;     //402pi/1024
   sin[202]  =  14'b11000011011111;     //404pi/1024
   cos[202]  =  14'b00010100110100;     //404pi/1024
   sin[203]  =  14'b11000011010111;     //406pi/1024
   cos[203]  =  14'b00010100011100;     //406pi/1024
   sin[204]  =  14'b11000011001111;     //408pi/1024
   cos[204]  =  14'b00010100000100;     //408pi/1024
   sin[205]  =  14'b11000011000111;     //410pi/1024
   cos[205]  =  14'b00010011101100;     //410pi/1024
   sin[206]  =  14'b11000010111111;     //412pi/1024
   cos[206]  =  14'b00010011010101;     //412pi/1024
   sin[207]  =  14'b11000010111000;     //414pi/1024
   cos[207]  =  14'b00010010111101;     //414pi/1024
   sin[208]  =  14'b11000010110000;     //416pi/1024
   cos[208]  =  14'b00010010100101;     //416pi/1024
   sin[209]  =  14'b11000010101001;     //418pi/1024
   cos[209]  =  14'b00010010001100;     //418pi/1024
   sin[210]  =  14'b11000010100010;     //420pi/1024
   cos[210]  =  14'b00010001110100;     //420pi/1024
   sin[211]  =  14'b11000010011011;     //422pi/1024
   cos[211]  =  14'b00010001011100;     //422pi/1024
   sin[212]  =  14'b11000010010100;     //424pi/1024
   cos[212]  =  14'b00010001000100;     //424pi/1024
   sin[213]  =  14'b11000010001110;     //426pi/1024
   cos[213]  =  14'b00010000101100;     //426pi/1024
   sin[214]  =  14'b11000010000111;     //428pi/1024
   cos[214]  =  14'b00010000010011;     //428pi/1024
   sin[215]  =  14'b11000010000001;     //430pi/1024
   cos[215]  =  14'b00001111111011;     //430pi/1024
   sin[216]  =  14'b11000001111011;     //432pi/1024
   cos[216]  =  14'b00001111100011;     //432pi/1024
   sin[217]  =  14'b11000001110101;     //434pi/1024
   cos[217]  =  14'b00001111001010;     //434pi/1024
   sin[218]  =  14'b11000001101111;     //436pi/1024
   cos[218]  =  14'b00001110110010;     //436pi/1024
   sin[219]  =  14'b11000001101001;     //438pi/1024
   cos[219]  =  14'b00001110011001;     //438pi/1024
   sin[220]  =  14'b11000001100100;     //440pi/1024
   cos[220]  =  14'b00001110000001;     //440pi/1024
   sin[221]  =  14'b11000001011110;     //442pi/1024
   cos[221]  =  14'b00001101101000;     //442pi/1024
   sin[222]  =  14'b11000001011001;     //444pi/1024
   cos[222]  =  14'b00001101010000;     //444pi/1024
   sin[223]  =  14'b11000001010100;     //446pi/1024
   cos[223]  =  14'b00001100110111;     //446pi/1024
   sin[224]  =  14'b11000001001111;     //448pi/1024
   cos[224]  =  14'b00001100011111;     //448pi/1024
   sin[225]  =  14'b11000001001010;     //450pi/1024
   cos[225]  =  14'b00001100000110;     //450pi/1024
   sin[226]  =  14'b11000001000101;     //452pi/1024
   cos[226]  =  14'b00001011101101;     //452pi/1024
   sin[227]  =  14'b11000001000001;     //454pi/1024
   cos[227]  =  14'b00001011010101;     //454pi/1024
   sin[228]  =  14'b11000000111100;     //456pi/1024
   cos[228]  =  14'b00001010111100;     //456pi/1024
   sin[229]  =  14'b11000000111000;     //458pi/1024
   cos[229]  =  14'b00001010100011;     //458pi/1024
   sin[230]  =  14'b11000000110100;     //460pi/1024
   cos[230]  =  14'b00001010001010;     //460pi/1024
   sin[231]  =  14'b11000000110000;     //462pi/1024
   cos[231]  =  14'b00001001110001;     //462pi/1024
   sin[232]  =  14'b11000000101100;     //464pi/1024
   cos[232]  =  14'b00001001011001;     //464pi/1024
   sin[233]  =  14'b11000000101001;     //466pi/1024
   cos[233]  =  14'b00001001000000;     //466pi/1024
   sin[234]  =  14'b11000000100101;     //468pi/1024
   cos[234]  =  14'b00001000100111;     //468pi/1024
   sin[235]  =  14'b11000000100010;     //470pi/1024
   cos[235]  =  14'b00001000001110;     //470pi/1024
   sin[236]  =  14'b11000000011111;     //472pi/1024
   cos[236]  =  14'b00000111110101;     //472pi/1024
   sin[237]  =  14'b11000000011100;     //474pi/1024
   cos[237]  =  14'b00000111011100;     //474pi/1024
   sin[238]  =  14'b11000000011001;     //476pi/1024
   cos[238]  =  14'b00000111000011;     //476pi/1024
   sin[239]  =  14'b11000000010110;     //478pi/1024
   cos[239]  =  14'b00000110101010;     //478pi/1024
   sin[240]  =  14'b11000000010100;     //480pi/1024
   cos[240]  =  14'b00000110010001;     //480pi/1024
   sin[241]  =  14'b11000000010001;     //482pi/1024
   cos[241]  =  14'b00000101111000;     //482pi/1024
   sin[242]  =  14'b11000000001111;     //484pi/1024
   cos[242]  =  14'b00000101011111;     //484pi/1024
   sin[243]  =  14'b11000000001101;     //486pi/1024
   cos[243]  =  14'b00000101000110;     //486pi/1024
   sin[244]  =  14'b11000000001011;     //488pi/1024
   cos[244]  =  14'b00000100101101;     //488pi/1024
   sin[245]  =  14'b11000000001001;     //490pi/1024
   cos[245]  =  14'b00000100010100;     //490pi/1024
   sin[246]  =  14'b11000000001000;     //492pi/1024
   cos[246]  =  14'b00000011111011;     //492pi/1024
   sin[247]  =  14'b11000000000110;     //494pi/1024
   cos[247]  =  14'b00000011100010;     //494pi/1024
   sin[248]  =  14'b11000000000101;     //496pi/1024
   cos[248]  =  14'b00000011001000;     //496pi/1024
   sin[249]  =  14'b11000000000100;     //498pi/1024
   cos[249]  =  14'b00000010101111;     //498pi/1024
   sin[250]  =  14'b11000000000011;     //500pi/1024
   cos[250]  =  14'b00000010010110;     //500pi/1024
   sin[251]  =  14'b11000000000010;     //502pi/1024
   cos[251]  =  14'b00000001111101;     //502pi/1024
   sin[252]  =  14'b11000000000001;     //504pi/1024
   cos[252]  =  14'b00000001100100;     //504pi/1024
   sin[253]  =  14'b11000000000001;     //506pi/1024
   cos[253]  =  14'b00000001001011;     //506pi/1024
   sin[254]  =  14'b11000000000000;     //508pi/1024
   cos[254]  =  14'b00000000110010;     //508pi/1024
   sin[255]  =  14'b11000000000000;     //510pi/1024
   cos[255]  =  14'b00000000011001;     //510pi/1024
   sin[256]  =  14'b11000000000000;     //512pi/1024
   cos[256]  =  14'b00000000000000;     //512pi/1024
   sin[257]  =  14'b11000000000000;     //514pi/1024
   cos[257]  =  14'b11111111100111;     //514pi/1024
   sin[258]  =  14'b11000000000000;     //516pi/1024
   cos[258]  =  14'b11111111001110;     //516pi/1024
   sin[259]  =  14'b11000000000001;     //518pi/1024
   cos[259]  =  14'b11111110110101;     //518pi/1024
   sin[260]  =  14'b11000000000001;     //520pi/1024
   cos[260]  =  14'b11111110011011;     //520pi/1024
   sin[261]  =  14'b11000000000010;     //522pi/1024
   cos[261]  =  14'b11111110000010;     //522pi/1024
   sin[262]  =  14'b11000000000011;     //524pi/1024
   cos[262]  =  14'b11111101101001;     //524pi/1024
   sin[263]  =  14'b11000000000100;     //526pi/1024
   cos[263]  =  14'b11111101010000;     //526pi/1024
   sin[264]  =  14'b11000000000101;     //528pi/1024
   cos[264]  =  14'b11111100110111;     //528pi/1024
   sin[265]  =  14'b11000000000110;     //530pi/1024
   cos[265]  =  14'b11111100011110;     //530pi/1024
   sin[266]  =  14'b11000000001000;     //532pi/1024
   cos[266]  =  14'b11111100000101;     //532pi/1024
   sin[267]  =  14'b11000000001001;     //534pi/1024
   cos[267]  =  14'b11111011101100;     //534pi/1024
   sin[268]  =  14'b11000000001011;     //536pi/1024
   cos[268]  =  14'b11111011010011;     //536pi/1024
   sin[269]  =  14'b11000000001101;     //538pi/1024
   cos[269]  =  14'b11111010111010;     //538pi/1024
   sin[270]  =  14'b11000000001111;     //540pi/1024
   cos[270]  =  14'b11111010100001;     //540pi/1024
   sin[271]  =  14'b11000000010001;     //542pi/1024
   cos[271]  =  14'b11111010001000;     //542pi/1024
   sin[272]  =  14'b11000000010100;     //544pi/1024
   cos[272]  =  14'b11111001101111;     //544pi/1024
   sin[273]  =  14'b11000000010110;     //546pi/1024
   cos[273]  =  14'b11111001010110;     //546pi/1024
   sin[274]  =  14'b11000000011001;     //548pi/1024
   cos[274]  =  14'b11111000111101;     //548pi/1024
   sin[275]  =  14'b11000000011100;     //550pi/1024
   cos[275]  =  14'b11111000100100;     //550pi/1024
   sin[276]  =  14'b11000000011111;     //552pi/1024
   cos[276]  =  14'b11111000001011;     //552pi/1024
   sin[277]  =  14'b11000000100010;     //554pi/1024
   cos[277]  =  14'b11110111110010;     //554pi/1024
   sin[278]  =  14'b11000000100101;     //556pi/1024
   cos[278]  =  14'b11110111011001;     //556pi/1024
   sin[279]  =  14'b11000000101001;     //558pi/1024
   cos[279]  =  14'b11110111000000;     //558pi/1024
   sin[280]  =  14'b11000000101100;     //560pi/1024
   cos[280]  =  14'b11110110100111;     //560pi/1024
   sin[281]  =  14'b11000000110000;     //562pi/1024
   cos[281]  =  14'b11110110001110;     //562pi/1024
   sin[282]  =  14'b11000000110100;     //564pi/1024
   cos[282]  =  14'b11110101110101;     //564pi/1024
   sin[283]  =  14'b11000000111000;     //566pi/1024
   cos[283]  =  14'b11110101011101;     //566pi/1024
   sin[284]  =  14'b11000000111100;     //568pi/1024
   cos[284]  =  14'b11110101000100;     //568pi/1024
   sin[285]  =  14'b11000001000001;     //570pi/1024
   cos[285]  =  14'b11110100101011;     //570pi/1024
   sin[286]  =  14'b11000001000101;     //572pi/1024
   cos[286]  =  14'b11110100010010;     //572pi/1024
   sin[287]  =  14'b11000001001010;     //574pi/1024
   cos[287]  =  14'b11110011111010;     //574pi/1024
   sin[288]  =  14'b11000001001111;     //576pi/1024
   cos[288]  =  14'b11110011100001;     //576pi/1024
   sin[289]  =  14'b11000001010100;     //578pi/1024
   cos[289]  =  14'b11110011001000;     //578pi/1024
   sin[290]  =  14'b11000001011001;     //580pi/1024
   cos[290]  =  14'b11110010110000;     //580pi/1024
   sin[291]  =  14'b11000001011110;     //582pi/1024
   cos[291]  =  14'b11110010010111;     //582pi/1024
   sin[292]  =  14'b11000001100100;     //584pi/1024
   cos[292]  =  14'b11110001111111;     //584pi/1024
   sin[293]  =  14'b11000001101001;     //586pi/1024
   cos[293]  =  14'b11110001100110;     //586pi/1024
   sin[294]  =  14'b11000001101111;     //588pi/1024
   cos[294]  =  14'b11110001001110;     //588pi/1024
   sin[295]  =  14'b11000001110101;     //590pi/1024
   cos[295]  =  14'b11110000110101;     //590pi/1024
   sin[296]  =  14'b11000001111011;     //592pi/1024
   cos[296]  =  14'b11110000011101;     //592pi/1024
   sin[297]  =  14'b11000010000001;     //594pi/1024
   cos[297]  =  14'b11110000000100;     //594pi/1024
   sin[298]  =  14'b11000010000111;     //596pi/1024
   cos[298]  =  14'b11101111101100;     //596pi/1024
   sin[299]  =  14'b11000010001110;     //598pi/1024
   cos[299]  =  14'b11101111010100;     //598pi/1024
   sin[300]  =  14'b11000010010100;     //600pi/1024
   cos[300]  =  14'b11101110111100;     //600pi/1024
   sin[301]  =  14'b11000010011011;     //602pi/1024
   cos[301]  =  14'b11101110100011;     //602pi/1024
   sin[302]  =  14'b11000010100010;     //604pi/1024
   cos[302]  =  14'b11101110001011;     //604pi/1024
   sin[303]  =  14'b11000010101001;     //606pi/1024
   cos[303]  =  14'b11101101110011;     //606pi/1024
   sin[304]  =  14'b11000010110000;     //608pi/1024
   cos[304]  =  14'b11101101011011;     //608pi/1024
   sin[305]  =  14'b11000010111000;     //610pi/1024
   cos[305]  =  14'b11101101000011;     //610pi/1024
   sin[306]  =  14'b11000010111111;     //612pi/1024
   cos[306]  =  14'b11101100101011;     //612pi/1024
   sin[307]  =  14'b11000011000111;     //614pi/1024
   cos[307]  =  14'b11101100010011;     //614pi/1024
   sin[308]  =  14'b11000011001111;     //616pi/1024
   cos[308]  =  14'b11101011111011;     //616pi/1024
   sin[309]  =  14'b11000011010111;     //618pi/1024
   cos[309]  =  14'b11101011100011;     //618pi/1024
   sin[310]  =  14'b11000011011111;     //620pi/1024
   cos[310]  =  14'b11101011001100;     //620pi/1024
   sin[311]  =  14'b11000011100111;     //622pi/1024
   cos[311]  =  14'b11101010110100;     //622pi/1024
   sin[312]  =  14'b11000011101111;     //624pi/1024
   cos[312]  =  14'b11101010011100;     //624pi/1024
   sin[313]  =  14'b11000011111000;     //626pi/1024
   cos[313]  =  14'b11101010000100;     //626pi/1024
   sin[314]  =  14'b11000100000001;     //628pi/1024
   cos[314]  =  14'b11101001101101;     //628pi/1024
   sin[315]  =  14'b11000100001001;     //630pi/1024
   cos[315]  =  14'b11101001010101;     //630pi/1024
   sin[316]  =  14'b11000100010010;     //632pi/1024
   cos[316]  =  14'b11101000111110;     //632pi/1024
   sin[317]  =  14'b11000100011100;     //634pi/1024
   cos[317]  =  14'b11101000100110;     //634pi/1024
   sin[318]  =  14'b11000100100101;     //636pi/1024
   cos[318]  =  14'b11101000001111;     //636pi/1024
   sin[319]  =  14'b11000100101110;     //638pi/1024
   cos[319]  =  14'b11100111111000;     //638pi/1024
   sin[320]  =  14'b11000100111000;     //640pi/1024
   cos[320]  =  14'b11100111100001;     //640pi/1024
   sin[321]  =  14'b11000101000001;     //642pi/1024
   cos[321]  =  14'b11100111001001;     //642pi/1024
   sin[322]  =  14'b11000101001011;     //644pi/1024
   cos[322]  =  14'b11100110110010;     //644pi/1024
   sin[323]  =  14'b11000101010101;     //646pi/1024
   cos[323]  =  14'b11100110011011;     //646pi/1024
   sin[324]  =  14'b11000101011111;     //648pi/1024
   cos[324]  =  14'b11100110000100;     //648pi/1024
   sin[325]  =  14'b11000101101010;     //650pi/1024
   cos[325]  =  14'b11100101101101;     //650pi/1024
   sin[326]  =  14'b11000101110100;     //652pi/1024
   cos[326]  =  14'b11100101010110;     //652pi/1024
   sin[327]  =  14'b11000101111111;     //654pi/1024
   cos[327]  =  14'b11100100111111;     //654pi/1024
   sin[328]  =  14'b11000110001001;     //656pi/1024
   cos[328]  =  14'b11100100101001;     //656pi/1024
   sin[329]  =  14'b11000110010100;     //658pi/1024
   cos[329]  =  14'b11100100010010;     //658pi/1024
   sin[330]  =  14'b11000110011111;     //660pi/1024
   cos[330]  =  14'b11100011111011;     //660pi/1024
   sin[331]  =  14'b11000110101010;     //662pi/1024
   cos[331]  =  14'b11100011100101;     //662pi/1024
   sin[332]  =  14'b11000110110101;     //664pi/1024
   cos[332]  =  14'b11100011001110;     //664pi/1024
   sin[333]  =  14'b11000111000001;     //666pi/1024
   cos[333]  =  14'b11100010111000;     //666pi/1024
   sin[334]  =  14'b11000111001100;     //668pi/1024
   cos[334]  =  14'b11100010100010;     //668pi/1024
   sin[335]  =  14'b11000111011000;     //670pi/1024
   cos[335]  =  14'b11100010001011;     //670pi/1024
   sin[336]  =  14'b11000111100100;     //672pi/1024
   cos[336]  =  14'b11100001110101;     //672pi/1024
   sin[337]  =  14'b11000111110000;     //674pi/1024
   cos[337]  =  14'b11100001011111;     //674pi/1024
   sin[338]  =  14'b11000111111100;     //676pi/1024
   cos[338]  =  14'b11100001001001;     //676pi/1024
   sin[339]  =  14'b11001000001000;     //678pi/1024
   cos[339]  =  14'b11100000110011;     //678pi/1024
   sin[340]  =  14'b11001000010100;     //680pi/1024
   cos[340]  =  14'b11100000011101;     //680pi/1024
   sin[341]  =  14'b11001000100001;     //682pi/1024
   cos[341]  =  14'b11100000000111;     //682pi/1024
   sin[342]  =  14'b11001000101101;     //684pi/1024
   cos[342]  =  14'b11011111110010;     //684pi/1024
   sin[343]  =  14'b11001000111010;     //686pi/1024
   cos[343]  =  14'b11011111011100;     //686pi/1024
   sin[344]  =  14'b11001001000111;     //688pi/1024
   cos[344]  =  14'b11011111000110;     //688pi/1024
   sin[345]  =  14'b11001001010100;     //690pi/1024
   cos[345]  =  14'b11011110110001;     //690pi/1024
   sin[346]  =  14'b11001001100001;     //692pi/1024
   cos[346]  =  14'b11011110011011;     //692pi/1024
   sin[347]  =  14'b11001001101110;     //694pi/1024
   cos[347]  =  14'b11011110000110;     //694pi/1024
   sin[348]  =  14'b11001001111011;     //696pi/1024
   cos[348]  =  14'b11011101110001;     //696pi/1024
   sin[349]  =  14'b11001010001001;     //698pi/1024
   cos[349]  =  14'b11011101011011;     //698pi/1024
   sin[350]  =  14'b11001010010111;     //700pi/1024
   cos[350]  =  14'b11011101000110;     //700pi/1024
   sin[351]  =  14'b11001010100100;     //702pi/1024
   cos[351]  =  14'b11011100110001;     //702pi/1024
   sin[352]  =  14'b11001010110010;     //704pi/1024
   cos[352]  =  14'b11011100011100;     //704pi/1024
   sin[353]  =  14'b11001011000000;     //706pi/1024
   cos[353]  =  14'b11011100001000;     //706pi/1024
   sin[354]  =  14'b11001011001110;     //708pi/1024
   cos[354]  =  14'b11011011110011;     //708pi/1024
   sin[355]  =  14'b11001011011101;     //710pi/1024
   cos[355]  =  14'b11011011011110;     //710pi/1024
   sin[356]  =  14'b11001011101011;     //712pi/1024
   cos[356]  =  14'b11011011001001;     //712pi/1024
   sin[357]  =  14'b11001011111010;     //714pi/1024
   cos[357]  =  14'b11011010110101;     //714pi/1024
   sin[358]  =  14'b11001100001000;     //716pi/1024
   cos[358]  =  14'b11011010100001;     //716pi/1024
   sin[359]  =  14'b11001100010111;     //718pi/1024
   cos[359]  =  14'b11011010001100;     //718pi/1024
   sin[360]  =  14'b11001100100110;     //720pi/1024
   cos[360]  =  14'b11011001111000;     //720pi/1024
   sin[361]  =  14'b11001100110101;     //722pi/1024
   cos[361]  =  14'b11011001100100;     //722pi/1024
   sin[362]  =  14'b11001101000100;     //724pi/1024
   cos[362]  =  14'b11011001010000;     //724pi/1024
   sin[363]  =  14'b11001101010100;     //726pi/1024
   cos[363]  =  14'b11011000111100;     //726pi/1024
   sin[364]  =  14'b11001101100011;     //728pi/1024
   cos[364]  =  14'b11011000101000;     //728pi/1024
   sin[365]  =  14'b11001101110010;     //730pi/1024
   cos[365]  =  14'b11011000010100;     //730pi/1024
   sin[366]  =  14'b11001110000010;     //732pi/1024
   cos[366]  =  14'b11011000000001;     //732pi/1024
   sin[367]  =  14'b11001110010010;     //734pi/1024
   cos[367]  =  14'b11010111101101;     //734pi/1024
   sin[368]  =  14'b11001110100010;     //736pi/1024
   cos[368]  =  14'b11010111011010;     //736pi/1024
   sin[369]  =  14'b11001110110010;     //738pi/1024
   cos[369]  =  14'b11010111000110;     //738pi/1024
   sin[370]  =  14'b11001111000010;     //740pi/1024
   cos[370]  =  14'b11010110110011;     //740pi/1024
   sin[371]  =  14'b11001111010010;     //742pi/1024
   cos[371]  =  14'b11010110100000;     //742pi/1024
   sin[372]  =  14'b11001111100010;     //744pi/1024
   cos[372]  =  14'b11010110001101;     //744pi/1024
   sin[373]  =  14'b11001111110011;     //746pi/1024
   cos[373]  =  14'b11010101111010;     //746pi/1024
   sin[374]  =  14'b11010000000100;     //748pi/1024
   cos[374]  =  14'b11010101100111;     //748pi/1024
   sin[375]  =  14'b11010000010100;     //750pi/1024
   cos[375]  =  14'b11010101010100;     //750pi/1024
   sin[376]  =  14'b11010000100101;     //752pi/1024
   cos[376]  =  14'b11010101000001;     //752pi/1024
   sin[377]  =  14'b11010000110110;     //754pi/1024
   cos[377]  =  14'b11010100101111;     //754pi/1024
   sin[378]  =  14'b11010001000111;     //756pi/1024
   cos[378]  =  14'b11010100011100;     //756pi/1024
   sin[379]  =  14'b11010001011000;     //758pi/1024
   cos[379]  =  14'b11010100001010;     //758pi/1024
   sin[380]  =  14'b11010001101001;     //760pi/1024
   cos[380]  =  14'b11010011111000;     //760pi/1024
   sin[381]  =  14'b11010001111011;     //762pi/1024
   cos[381]  =  14'b11010011100101;     //762pi/1024
   sin[382]  =  14'b11010010001100;     //764pi/1024
   cos[382]  =  14'b11010011010011;     //764pi/1024
   sin[383]  =  14'b11010010011110;     //766pi/1024
   cos[383]  =  14'b11010011000010;     //766pi/1024
   sin[384]  =  14'b11010010110000;     //768pi/1024
   cos[384]  =  14'b11010010110000;     //768pi/1024
   sin[385]  =  14'b11010011000010;     //770pi/1024
   cos[385]  =  14'b11010010011110;     //770pi/1024
   sin[386]  =  14'b11010011010011;     //772pi/1024
   cos[386]  =  14'b11010010001100;     //772pi/1024
   sin[387]  =  14'b11010011100101;     //774pi/1024
   cos[387]  =  14'b11010001111011;     //774pi/1024
   sin[388]  =  14'b11010011111000;     //776pi/1024
   cos[388]  =  14'b11010001101001;     //776pi/1024
   sin[389]  =  14'b11010100001010;     //778pi/1024
   cos[389]  =  14'b11010001011000;     //778pi/1024
   sin[390]  =  14'b11010100011100;     //780pi/1024
   cos[390]  =  14'b11010001000111;     //780pi/1024
   sin[391]  =  14'b11010100101111;     //782pi/1024
   cos[391]  =  14'b11010000110110;     //782pi/1024
   sin[392]  =  14'b11010101000001;     //784pi/1024
   cos[392]  =  14'b11010000100101;     //784pi/1024
   sin[393]  =  14'b11010101010100;     //786pi/1024
   cos[393]  =  14'b11010000010100;     //786pi/1024
   sin[394]  =  14'b11010101100111;     //788pi/1024
   cos[394]  =  14'b11010000000100;     //788pi/1024
   sin[395]  =  14'b11010101111010;     //790pi/1024
   cos[395]  =  14'b11001111110011;     //790pi/1024
   sin[396]  =  14'b11010110001101;     //792pi/1024
   cos[396]  =  14'b11001111100010;     //792pi/1024
   sin[397]  =  14'b11010110100000;     //794pi/1024
   cos[397]  =  14'b11001111010010;     //794pi/1024
   sin[398]  =  14'b11010110110011;     //796pi/1024
   cos[398]  =  14'b11001111000010;     //796pi/1024
   sin[399]  =  14'b11010111000110;     //798pi/1024
   cos[399]  =  14'b11001110110010;     //798pi/1024
   sin[400]  =  14'b11010111011010;     //800pi/1024
   cos[400]  =  14'b11001110100010;     //800pi/1024
   sin[401]  =  14'b11010111101101;     //802pi/1024
   cos[401]  =  14'b11001110010010;     //802pi/1024
   sin[402]  =  14'b11011000000001;     //804pi/1024
   cos[402]  =  14'b11001110000010;     //804pi/1024
   sin[403]  =  14'b11011000010100;     //806pi/1024
   cos[403]  =  14'b11001101110010;     //806pi/1024
   sin[404]  =  14'b11011000101000;     //808pi/1024
   cos[404]  =  14'b11001101100011;     //808pi/1024
   sin[405]  =  14'b11011000111100;     //810pi/1024
   cos[405]  =  14'b11001101010100;     //810pi/1024
   sin[406]  =  14'b11011001010000;     //812pi/1024
   cos[406]  =  14'b11001101000100;     //812pi/1024
   sin[407]  =  14'b11011001100100;     //814pi/1024
   cos[407]  =  14'b11001100110101;     //814pi/1024
   sin[408]  =  14'b11011001111000;     //816pi/1024
   cos[408]  =  14'b11001100100110;     //816pi/1024
   sin[409]  =  14'b11011010001100;     //818pi/1024
   cos[409]  =  14'b11001100010111;     //818pi/1024
   sin[410]  =  14'b11011010100001;     //820pi/1024
   cos[410]  =  14'b11001100001000;     //820pi/1024
   sin[411]  =  14'b11011010110101;     //822pi/1024
   cos[411]  =  14'b11001011111010;     //822pi/1024
   sin[412]  =  14'b11011011001001;     //824pi/1024
   cos[412]  =  14'b11001011101011;     //824pi/1024
   sin[413]  =  14'b11011011011110;     //826pi/1024
   cos[413]  =  14'b11001011011101;     //826pi/1024
   sin[414]  =  14'b11011011110011;     //828pi/1024
   cos[414]  =  14'b11001011001110;     //828pi/1024
   sin[415]  =  14'b11011100001000;     //830pi/1024
   cos[415]  =  14'b11001011000000;     //830pi/1024
   sin[416]  =  14'b11011100011100;     //832pi/1024
   cos[416]  =  14'b11001010110010;     //832pi/1024
   sin[417]  =  14'b11011100110001;     //834pi/1024
   cos[417]  =  14'b11001010100100;     //834pi/1024
   sin[418]  =  14'b11011101000110;     //836pi/1024
   cos[418]  =  14'b11001010010111;     //836pi/1024
   sin[419]  =  14'b11011101011011;     //838pi/1024
   cos[419]  =  14'b11001010001001;     //838pi/1024
   sin[420]  =  14'b11011101110001;     //840pi/1024
   cos[420]  =  14'b11001001111011;     //840pi/1024
   sin[421]  =  14'b11011110000110;     //842pi/1024
   cos[421]  =  14'b11001001101110;     //842pi/1024
   sin[422]  =  14'b11011110011011;     //844pi/1024
   cos[422]  =  14'b11001001100001;     //844pi/1024
   sin[423]  =  14'b11011110110001;     //846pi/1024
   cos[423]  =  14'b11001001010100;     //846pi/1024
   sin[424]  =  14'b11011111000110;     //848pi/1024
   cos[424]  =  14'b11001001000111;     //848pi/1024
   sin[425]  =  14'b11011111011100;     //850pi/1024
   cos[425]  =  14'b11001000111010;     //850pi/1024
   sin[426]  =  14'b11011111110010;     //852pi/1024
   cos[426]  =  14'b11001000101101;     //852pi/1024
   sin[427]  =  14'b11100000000111;     //854pi/1024
   cos[427]  =  14'b11001000100001;     //854pi/1024
   sin[428]  =  14'b11100000011101;     //856pi/1024
   cos[428]  =  14'b11001000010100;     //856pi/1024
   sin[429]  =  14'b11100000110011;     //858pi/1024
   cos[429]  =  14'b11001000001000;     //858pi/1024
   sin[430]  =  14'b11100001001001;     //860pi/1024
   cos[430]  =  14'b11000111111100;     //860pi/1024
   sin[431]  =  14'b11100001011111;     //862pi/1024
   cos[431]  =  14'b11000111110000;     //862pi/1024
   sin[432]  =  14'b11100001110101;     //864pi/1024
   cos[432]  =  14'b11000111100100;     //864pi/1024
   sin[433]  =  14'b11100010001011;     //866pi/1024
   cos[433]  =  14'b11000111011000;     //866pi/1024
   sin[434]  =  14'b11100010100010;     //868pi/1024
   cos[434]  =  14'b11000111001100;     //868pi/1024
   sin[435]  =  14'b11100010111000;     //870pi/1024
   cos[435]  =  14'b11000111000001;     //870pi/1024
   sin[436]  =  14'b11100011001110;     //872pi/1024
   cos[436]  =  14'b11000110110101;     //872pi/1024
   sin[437]  =  14'b11100011100101;     //874pi/1024
   cos[437]  =  14'b11000110101010;     //874pi/1024
   sin[438]  =  14'b11100011111011;     //876pi/1024
   cos[438]  =  14'b11000110011111;     //876pi/1024
   sin[439]  =  14'b11100100010010;     //878pi/1024
   cos[439]  =  14'b11000110010100;     //878pi/1024
   sin[440]  =  14'b11100100101001;     //880pi/1024
   cos[440]  =  14'b11000110001001;     //880pi/1024
   sin[441]  =  14'b11100100111111;     //882pi/1024
   cos[441]  =  14'b11000101111111;     //882pi/1024
   sin[442]  =  14'b11100101010110;     //884pi/1024
   cos[442]  =  14'b11000101110100;     //884pi/1024
   sin[443]  =  14'b11100101101101;     //886pi/1024
   cos[443]  =  14'b11000101101010;     //886pi/1024
   sin[444]  =  14'b11100110000100;     //888pi/1024
   cos[444]  =  14'b11000101011111;     //888pi/1024
   sin[445]  =  14'b11100110011011;     //890pi/1024
   cos[445]  =  14'b11000101010101;     //890pi/1024
   sin[446]  =  14'b11100110110010;     //892pi/1024
   cos[446]  =  14'b11000101001011;     //892pi/1024
   sin[447]  =  14'b11100111001001;     //894pi/1024
   cos[447]  =  14'b11000101000001;     //894pi/1024
   sin[448]  =  14'b11100111100001;     //896pi/1024
   cos[448]  =  14'b11000100111000;     //896pi/1024
   sin[449]  =  14'b11100111111000;     //898pi/1024
   cos[449]  =  14'b11000100101110;     //898pi/1024
   sin[450]  =  14'b11101000001111;     //900pi/1024
   cos[450]  =  14'b11000100100101;     //900pi/1024
   sin[451]  =  14'b11101000100110;     //902pi/1024
   cos[451]  =  14'b11000100011100;     //902pi/1024
   sin[452]  =  14'b11101000111110;     //904pi/1024
   cos[452]  =  14'b11000100010010;     //904pi/1024
   sin[453]  =  14'b11101001010101;     //906pi/1024
   cos[453]  =  14'b11000100001001;     //906pi/1024
   sin[454]  =  14'b11101001101101;     //908pi/1024
   cos[454]  =  14'b11000100000001;     //908pi/1024
   sin[455]  =  14'b11101010000100;     //910pi/1024
   cos[455]  =  14'b11000011111000;     //910pi/1024
   sin[456]  =  14'b11101010011100;     //912pi/1024
   cos[456]  =  14'b11000011101111;     //912pi/1024
   sin[457]  =  14'b11101010110100;     //914pi/1024
   cos[457]  =  14'b11000011100111;     //914pi/1024
   sin[458]  =  14'b11101011001100;     //916pi/1024
   cos[458]  =  14'b11000011011111;     //916pi/1024
   sin[459]  =  14'b11101011100011;     //918pi/1024
   cos[459]  =  14'b11000011010111;     //918pi/1024
   sin[460]  =  14'b11101011111011;     //920pi/1024
   cos[460]  =  14'b11000011001111;     //920pi/1024
   sin[461]  =  14'b11101100010011;     //922pi/1024
   cos[461]  =  14'b11000011000111;     //922pi/1024
   sin[462]  =  14'b11101100101011;     //924pi/1024
   cos[462]  =  14'b11000010111111;     //924pi/1024
   sin[463]  =  14'b11101101000011;     //926pi/1024
   cos[463]  =  14'b11000010111000;     //926pi/1024
   sin[464]  =  14'b11101101011011;     //928pi/1024
   cos[464]  =  14'b11000010110000;     //928pi/1024
   sin[465]  =  14'b11101101110011;     //930pi/1024
   cos[465]  =  14'b11000010101001;     //930pi/1024
   sin[466]  =  14'b11101110001011;     //932pi/1024
   cos[466]  =  14'b11000010100010;     //932pi/1024
   sin[467]  =  14'b11101110100011;     //934pi/1024
   cos[467]  =  14'b11000010011011;     //934pi/1024
   sin[468]  =  14'b11101110111100;     //936pi/1024
   cos[468]  =  14'b11000010010100;     //936pi/1024
   sin[469]  =  14'b11101111010100;     //938pi/1024
   cos[469]  =  14'b11000010001110;     //938pi/1024
   sin[470]  =  14'b11101111101100;     //940pi/1024
   cos[470]  =  14'b11000010000111;     //940pi/1024
   sin[471]  =  14'b11110000000100;     //942pi/1024
   cos[471]  =  14'b11000010000001;     //942pi/1024
   sin[472]  =  14'b11110000011101;     //944pi/1024
   cos[472]  =  14'b11000001111011;     //944pi/1024
   sin[473]  =  14'b11110000110101;     //946pi/1024
   cos[473]  =  14'b11000001110101;     //946pi/1024
   sin[474]  =  14'b11110001001110;     //948pi/1024
   cos[474]  =  14'b11000001101111;     //948pi/1024
   sin[475]  =  14'b11110001100110;     //950pi/1024
   cos[475]  =  14'b11000001101001;     //950pi/1024
   sin[476]  =  14'b11110001111111;     //952pi/1024
   cos[476]  =  14'b11000001100100;     //952pi/1024
   sin[477]  =  14'b11110010010111;     //954pi/1024
   cos[477]  =  14'b11000001011110;     //954pi/1024
   sin[478]  =  14'b11110010110000;     //956pi/1024
   cos[478]  =  14'b11000001011001;     //956pi/1024
   sin[479]  =  14'b11110011001000;     //958pi/1024
   cos[479]  =  14'b11000001010100;     //958pi/1024
   sin[480]  =  14'b11110011100001;     //960pi/1024
   cos[480]  =  14'b11000001001111;     //960pi/1024
   sin[481]  =  14'b11110011111010;     //962pi/1024
   cos[481]  =  14'b11000001001010;     //962pi/1024
   sin[482]  =  14'b11110100010010;     //964pi/1024
   cos[482]  =  14'b11000001000101;     //964pi/1024
   sin[483]  =  14'b11110100101011;     //966pi/1024
   cos[483]  =  14'b11000001000001;     //966pi/1024
   sin[484]  =  14'b11110101000100;     //968pi/1024
   cos[484]  =  14'b11000000111100;     //968pi/1024
   sin[485]  =  14'b11110101011101;     //970pi/1024
   cos[485]  =  14'b11000000111000;     //970pi/1024
   sin[486]  =  14'b11110101110101;     //972pi/1024
   cos[486]  =  14'b11000000110100;     //972pi/1024
   sin[487]  =  14'b11110110001110;     //974pi/1024
   cos[487]  =  14'b11000000110000;     //974pi/1024
   sin[488]  =  14'b11110110100111;     //976pi/1024
   cos[488]  =  14'b11000000101100;     //976pi/1024
   sin[489]  =  14'b11110111000000;     //978pi/1024
   cos[489]  =  14'b11000000101001;     //978pi/1024
   sin[490]  =  14'b11110111011001;     //980pi/1024
   cos[490]  =  14'b11000000100101;     //980pi/1024
   sin[491]  =  14'b11110111110010;     //982pi/1024
   cos[491]  =  14'b11000000100010;     //982pi/1024
   sin[492]  =  14'b11111000001011;     //984pi/1024
   cos[492]  =  14'b11000000011111;     //984pi/1024
   sin[493]  =  14'b11111000100100;     //986pi/1024
   cos[493]  =  14'b11000000011100;     //986pi/1024
   sin[494]  =  14'b11111000111101;     //988pi/1024
   cos[494]  =  14'b11000000011001;     //988pi/1024
   sin[495]  =  14'b11111001010110;     //990pi/1024
   cos[495]  =  14'b11000000010110;     //990pi/1024
   sin[496]  =  14'b11111001101111;     //992pi/1024
   cos[496]  =  14'b11000000010100;     //992pi/1024
   sin[497]  =  14'b11111010001000;     //994pi/1024
   cos[497]  =  14'b11000000010001;     //994pi/1024
   sin[498]  =  14'b11111010100001;     //996pi/1024
   cos[498]  =  14'b11000000001111;     //996pi/1024
   sin[499]  =  14'b11111010111010;     //998pi/1024
   cos[499]  =  14'b11000000001101;     //998pi/1024
   sin[500]  =  14'b11111011010011;     //1000pi/1024
   cos[500]  =  14'b11000000001011;     //1000pi/1024
   sin[501]  =  14'b11111011101100;     //1002pi/1024
   cos[501]  =  14'b11000000001001;     //1002pi/1024
   sin[502]  =  14'b11111100000101;     //1004pi/1024
   cos[502]  =  14'b11000000001000;     //1004pi/1024
   sin[503]  =  14'b11111100011110;     //1006pi/1024
   cos[503]  =  14'b11000000000110;     //1006pi/1024
   sin[504]  =  14'b11111100110111;     //1008pi/1024
   cos[504]  =  14'b11000000000101;     //1008pi/1024
   sin[505]  =  14'b11111101010000;     //1010pi/1024
   cos[505]  =  14'b11000000000100;     //1010pi/1024
   sin[506]  =  14'b11111101101001;     //1012pi/1024
   cos[506]  =  14'b11000000000011;     //1012pi/1024
   sin[507]  =  14'b11111110000010;     //1014pi/1024
   cos[507]  =  14'b11000000000010;     //1014pi/1024
   sin[508]  =  14'b11111110011011;     //1016pi/1024
   cos[508]  =  14'b11000000000001;     //1016pi/1024
   sin[509]  =  14'b11111110110101;     //1018pi/1024
   cos[509]  =  14'b11000000000001;     //1018pi/1024
   sin[510]  =  14'b11111111001110;     //1020pi/1024
   cos[510]  =  14'b11000000000000;     //1020pi/1024
   sin[511]  =  14'b11111111100111;     //1022pi/1024
   cos[511]  =  14'b11000000000000;     //1022pi/1024
end
endmodule