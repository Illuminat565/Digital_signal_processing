module  M_TWIDLE_0_05_v #(parameter stage_FFT = 2, SIZE =10, word_length_tw = 14) (
    input            clk,
    input            en_rd, 
    input   [stage_FFT-2:0]   rd_ptr_angle,

    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );



reg signed [word_length_tw-1:0]  m_cos  [511:0];
reg signed [word_length_tw-1:0]  m_sin  [511:0];


//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd ) begin
                  cos_data           <= m_cos   [rd_ptr_angle];
                  sin_data           <= m_sin   [rd_ptr_angle];
             end 
        end

//----------------------------------------------------------------------------------------
initial begin

   m_sin[0]  =  14'b00000000000000;     //0pi/512
   m_cos[0]  =  14'b01000000000000;     //0pi/512
   m_sin[1]  =  14'b11111111101000;     //1pi/512
   m_cos[1]  =  14'b00111111111111;     //1pi/512
   m_sin[2]  =  14'b11111111010000;     //2pi/512
   m_cos[2]  =  14'b00111111111111;     //2pi/512
   m_sin[3]  =  14'b11111110111000;     //3pi/512
   m_cos[3]  =  14'b00111111111111;     //3pi/512
   m_sin[4]  =  14'b11111110100001;     //4pi/512
   m_cos[4]  =  14'b00111111111110;     //4pi/512
   m_sin[5]  =  14'b11111110001001;     //5pi/512
   m_cos[5]  =  14'b00111111111110;     //5pi/512
   m_sin[6]  =  14'b11111101110001;     //6pi/512
   m_cos[6]  =  14'b00111111111101;     //6pi/512
   m_sin[7]  =  14'b11111101011001;     //7pi/512
   m_cos[7]  =  14'b00111111111100;     //7pi/512
   m_sin[8]  =  14'b11111101000001;     //8pi/512
   m_cos[8]  =  14'b00111111111011;     //8pi/512
   m_sin[9]  =  14'b11111100101001;     //9pi/512
   m_cos[9]  =  14'b00111111111010;     //9pi/512
   m_sin[10]  =  14'b11111100010001;     //10pi/512
   m_cos[10]  =  14'b00111111111001;     //10pi/512
   m_sin[11]  =  14'b11111011111010;     //11pi/512
   m_cos[11]  =  14'b00111111110111;     //11pi/512
   m_sin[12]  =  14'b11111011100010;     //12pi/512
   m_cos[12]  =  14'b00111111110101;     //12pi/512
   m_sin[13]  =  14'b11111011001010;     //13pi/512
   m_cos[13]  =  14'b00111111110100;     //13pi/512
   m_sin[14]  =  14'b11111010110010;     //14pi/512
   m_cos[14]  =  14'b00111111110010;     //14pi/512
   m_sin[15]  =  14'b11111010011010;     //15pi/512
   m_cos[15]  =  14'b00111111110000;     //15pi/512
   m_sin[16]  =  14'b11111010000011;     //16pi/512
   m_cos[16]  =  14'b00111111101110;     //16pi/512
   m_sin[17]  =  14'b11111001101011;     //17pi/512
   m_cos[17]  =  14'b00111111101011;     //17pi/512
   m_sin[18]  =  14'b11111001010011;     //18pi/512
   m_cos[18]  =  14'b00111111101001;     //18pi/512
   m_sin[19]  =  14'b11111000111011;     //19pi/512
   m_cos[19]  =  14'b00111111100110;     //19pi/512
   m_sin[20]  =  14'b11111000100100;     //20pi/512
   m_cos[20]  =  14'b00111111100100;     //20pi/512
   m_sin[21]  =  14'b11111000001100;     //21pi/512
   m_cos[21]  =  14'b00111111100001;     //21pi/512
   m_sin[22]  =  14'b11110111110100;     //22pi/512
   m_cos[22]  =  14'b00111111011110;     //22pi/512
   m_sin[23]  =  14'b11110111011100;     //23pi/512
   m_cos[23]  =  14'b00111111011011;     //23pi/512
   m_sin[24]  =  14'b11110111000101;     //24pi/512
   m_cos[24]  =  14'b00111111010111;     //24pi/512
   m_sin[25]  =  14'b11110110101101;     //25pi/512
   m_cos[25]  =  14'b00111111010100;     //25pi/512
   m_sin[26]  =  14'b11110110010110;     //26pi/512
   m_cos[26]  =  14'b00111111010001;     //26pi/512
   m_sin[27]  =  14'b11110101111110;     //27pi/512
   m_cos[27]  =  14'b00111111001101;     //27pi/512
   m_sin[28]  =  14'b11110101100110;     //28pi/512
   m_cos[28]  =  14'b00111111001001;     //28pi/512
   m_sin[29]  =  14'b11110101001111;     //29pi/512
   m_cos[29]  =  14'b00111111000101;     //29pi/512
   m_sin[30]  =  14'b11110100110111;     //30pi/512
   m_cos[30]  =  14'b00111111000001;     //30pi/512
   m_sin[31]  =  14'b11110100100000;     //31pi/512
   m_cos[31]  =  14'b00111110111101;     //31pi/512
   m_sin[32]  =  14'b11110100001000;     //32pi/512
   m_cos[32]  =  14'b00111110111000;     //32pi/512
   m_sin[33]  =  14'b11110011110001;     //33pi/512
   m_cos[33]  =  14'b00111110110100;     //33pi/512
   m_sin[34]  =  14'b11110011011010;     //34pi/512
   m_cos[34]  =  14'b00111110101111;     //34pi/512
   m_sin[35]  =  14'b11110011000010;     //35pi/512
   m_cos[35]  =  14'b00111110101011;     //35pi/512
   m_sin[36]  =  14'b11110010101011;     //36pi/512
   m_cos[36]  =  14'b00111110100110;     //36pi/512
   m_sin[37]  =  14'b11110010010011;     //37pi/512
   m_cos[37]  =  14'b00111110100001;     //37pi/512
   m_sin[38]  =  14'b11110001111100;     //38pi/512
   m_cos[38]  =  14'b00111110011011;     //38pi/512
   m_sin[39]  =  14'b11110001100101;     //39pi/512
   m_cos[39]  =  14'b00111110010110;     //39pi/512
   m_sin[40]  =  14'b11110001001110;     //40pi/512
   m_cos[40]  =  14'b00111110010001;     //40pi/512
   m_sin[41]  =  14'b11110000110110;     //41pi/512
   m_cos[41]  =  14'b00111110001011;     //41pi/512
   m_sin[42]  =  14'b11110000011111;     //42pi/512
   m_cos[42]  =  14'b00111110000101;     //42pi/512
   m_sin[43]  =  14'b11110000001000;     //43pi/512
   m_cos[43]  =  14'b00111110000000;     //43pi/512
   m_sin[44]  =  14'b11101111110001;     //44pi/512
   m_cos[44]  =  14'b00111101111010;     //44pi/512
   m_sin[45]  =  14'b11101111011010;     //45pi/512
   m_cos[45]  =  14'b00111101110011;     //45pi/512
   m_sin[46]  =  14'b11101111000011;     //46pi/512
   m_cos[46]  =  14'b00111101101101;     //46pi/512
   m_sin[47]  =  14'b11101110101100;     //47pi/512
   m_cos[47]  =  14'b00111101100111;     //47pi/512
   m_sin[48]  =  14'b11101110010101;     //48pi/512
   m_cos[48]  =  14'b00111101100000;     //48pi/512
   m_sin[49]  =  14'b11101101111110;     //49pi/512
   m_cos[49]  =  14'b00111101011010;     //49pi/512
   m_sin[50]  =  14'b11101101100111;     //50pi/512
   m_cos[50]  =  14'b00111101010011;     //50pi/512
   m_sin[51]  =  14'b11101101010000;     //51pi/512
   m_cos[51]  =  14'b00111101001100;     //51pi/512
   m_sin[52]  =  14'b11101100111001;     //52pi/512
   m_cos[52]  =  14'b00111101000101;     //52pi/512
   m_sin[53]  =  14'b11101100100011;     //53pi/512
   m_cos[53]  =  14'b00111100111110;     //53pi/512
   m_sin[54]  =  14'b11101100001100;     //54pi/512
   m_cos[54]  =  14'b00111100110110;     //54pi/512
   m_sin[55]  =  14'b11101011110101;     //55pi/512
   m_cos[55]  =  14'b00111100101111;     //55pi/512
   m_sin[56]  =  14'b11101011011111;     //56pi/512
   m_cos[56]  =  14'b00111100100111;     //56pi/512
   m_sin[57]  =  14'b11101011001000;     //57pi/512
   m_cos[57]  =  14'b00111100011111;     //57pi/512
   m_sin[58]  =  14'b11101010110001;     //58pi/512
   m_cos[58]  =  14'b00111100011000;     //58pi/512
   m_sin[59]  =  14'b11101010011011;     //59pi/512
   m_cos[59]  =  14'b00111100010000;     //59pi/512
   m_sin[60]  =  14'b11101010000100;     //60pi/512
   m_cos[60]  =  14'b00111100001000;     //60pi/512
   m_sin[61]  =  14'b11101001101110;     //61pi/512
   m_cos[61]  =  14'b00111011111111;     //61pi/512
   m_sin[62]  =  14'b11101001011000;     //62pi/512
   m_cos[62]  =  14'b00111011110111;     //62pi/512
   m_sin[63]  =  14'b11101001000001;     //63pi/512
   m_cos[63]  =  14'b00111011101110;     //63pi/512
   m_sin[64]  =  14'b11101000101011;     //64pi/512
   m_cos[64]  =  14'b00111011100110;     //64pi/512
   m_sin[65]  =  14'b11101000010101;     //65pi/512
   m_cos[65]  =  14'b00111011011101;     //65pi/512
   m_sin[66]  =  14'b11100111111111;     //66pi/512
   m_cos[66]  =  14'b00111011010100;     //66pi/512
   m_sin[67]  =  14'b11100111101001;     //67pi/512
   m_cos[67]  =  14'b00111011001011;     //67pi/512
   m_sin[68]  =  14'b11100111010011;     //68pi/512
   m_cos[68]  =  14'b00111011000010;     //68pi/512
   m_sin[69]  =  14'b11100110111101;     //69pi/512
   m_cos[69]  =  14'b00111010111001;     //69pi/512
   m_sin[70]  =  14'b11100110100111;     //70pi/512
   m_cos[70]  =  14'b00111010101111;     //70pi/512
   m_sin[71]  =  14'b11100110010001;     //71pi/512
   m_cos[71]  =  14'b00111010100110;     //71pi/512
   m_sin[72]  =  14'b11100101111011;     //72pi/512
   m_cos[72]  =  14'b00111010011100;     //72pi/512
   m_sin[73]  =  14'b11100101100101;     //73pi/512
   m_cos[73]  =  14'b00111010010010;     //73pi/512
   m_sin[74]  =  14'b11100101001111;     //74pi/512
   m_cos[74]  =  14'b00111010001000;     //74pi/512
   m_sin[75]  =  14'b11100100111010;     //75pi/512
   m_cos[75]  =  14'b00111001111110;     //75pi/512
   m_sin[76]  =  14'b11100100100100;     //76pi/512
   m_cos[76]  =  14'b00111001110100;     //76pi/512
   m_sin[77]  =  14'b11100100001111;     //77pi/512
   m_cos[77]  =  14'b00111001101010;     //77pi/512
   m_sin[78]  =  14'b11100011111001;     //78pi/512
   m_cos[78]  =  14'b00111001011111;     //78pi/512
   m_sin[79]  =  14'b11100011100100;     //79pi/512
   m_cos[79]  =  14'b00111001010101;     //79pi/512
   m_sin[80]  =  14'b11100011001110;     //80pi/512
   m_cos[80]  =  14'b00111001001010;     //80pi/512
   m_sin[81]  =  14'b11100010111001;     //81pi/512
   m_cos[81]  =  14'b00111000111111;     //81pi/512
   m_sin[82]  =  14'b11100010100100;     //82pi/512
   m_cos[82]  =  14'b00111000110100;     //82pi/512
   m_sin[83]  =  14'b11100010001111;     //83pi/512
   m_cos[83]  =  14'b00111000101001;     //83pi/512
   m_sin[84]  =  14'b11100001111010;     //84pi/512
   m_cos[84]  =  14'b00111000011110;     //84pi/512
   m_sin[85]  =  14'b11100001100101;     //85pi/512
   m_cos[85]  =  14'b00111000010011;     //85pi/512
   m_sin[86]  =  14'b11100001010000;     //86pi/512
   m_cos[86]  =  14'b00111000001000;     //86pi/512
   m_sin[87]  =  14'b11100000111011;     //87pi/512
   m_cos[87]  =  14'b00110111111100;     //87pi/512
   m_sin[88]  =  14'b11100000100110;     //88pi/512
   m_cos[88]  =  14'b00110111110000;     //88pi/512
   m_sin[89]  =  14'b11100000010001;     //89pi/512
   m_cos[89]  =  14'b00110111100101;     //89pi/512
   m_sin[90]  =  14'b11011111111100;     //90pi/512
   m_cos[90]  =  14'b00110111011001;     //90pi/512
   m_sin[91]  =  14'b11011111101000;     //91pi/512
   m_cos[91]  =  14'b00110111001101;     //91pi/512
   m_sin[92]  =  14'b11011111010011;     //92pi/512
   m_cos[92]  =  14'b00110111000000;     //92pi/512
   m_sin[93]  =  14'b11011110111111;     //93pi/512
   m_cos[93]  =  14'b00110110110100;     //93pi/512
   m_sin[94]  =  14'b11011110101010;     //94pi/512
   m_cos[94]  =  14'b00110110101000;     //94pi/512
   m_sin[95]  =  14'b11011110010110;     //95pi/512
   m_cos[95]  =  14'b00110110011011;     //95pi/512
   m_sin[96]  =  14'b11011110000010;     //96pi/512
   m_cos[96]  =  14'b00110110001111;     //96pi/512
   m_sin[97]  =  14'b11011101101101;     //97pi/512
   m_cos[97]  =  14'b00110110000010;     //97pi/512
   m_sin[98]  =  14'b11011101011001;     //98pi/512
   m_cos[98]  =  14'b00110101110101;     //98pi/512
   m_sin[99]  =  14'b11011101000101;     //99pi/512
   m_cos[99]  =  14'b00110101101000;     //99pi/512
   m_sin[100]  =  14'b11011100110001;     //100pi/512
   m_cos[100]  =  14'b00110101011011;     //100pi/512
   m_sin[101]  =  14'b11011100011101;     //101pi/512
   m_cos[101]  =  14'b00110101001110;     //101pi/512
   m_sin[102]  =  14'b11011100001010;     //102pi/512
   m_cos[102]  =  14'b00110101000001;     //102pi/512
   m_sin[103]  =  14'b11011011110110;     //103pi/512
   m_cos[103]  =  14'b00110100110011;     //103pi/512
   m_sin[104]  =  14'b11011011100010;     //104pi/512
   m_cos[104]  =  14'b00110100100110;     //104pi/512
   m_sin[105]  =  14'b11011011001111;     //105pi/512
   m_cos[105]  =  14'b00110100011000;     //105pi/512
   m_sin[106]  =  14'b11011010111011;     //106pi/512
   m_cos[106]  =  14'b00110100001010;     //106pi/512
   m_sin[107]  =  14'b11011010101000;     //107pi/512
   m_cos[107]  =  14'b00110011111100;     //107pi/512
   m_sin[108]  =  14'b11011010010100;     //108pi/512
   m_cos[108]  =  14'b00110011101110;     //108pi/512
   m_sin[109]  =  14'b11011010000001;     //109pi/512
   m_cos[109]  =  14'b00110011100000;     //109pi/512
   m_sin[110]  =  14'b11011001101110;     //110pi/512
   m_cos[110]  =  14'b00110011010010;     //110pi/512
   m_sin[111]  =  14'b11011001011011;     //111pi/512
   m_cos[111]  =  14'b00110011000100;     //111pi/512
   m_sin[112]  =  14'b11011001001000;     //112pi/512
   m_cos[112]  =  14'b00110010110101;     //112pi/512
   m_sin[113]  =  14'b11011000110101;     //113pi/512
   m_cos[113]  =  14'b00110010100111;     //113pi/512
   m_sin[114]  =  14'b11011000100010;     //114pi/512
   m_cos[114]  =  14'b00110010011000;     //114pi/512
   m_sin[115]  =  14'b11011000001111;     //115pi/512
   m_cos[115]  =  14'b00110010001001;     //115pi/512
   m_sin[116]  =  14'b11010111111101;     //116pi/512
   m_cos[116]  =  14'b00110001111010;     //116pi/512
   m_sin[117]  =  14'b11010111101010;     //117pi/512
   m_cos[117]  =  14'b00110001101011;     //117pi/512
   m_sin[118]  =  14'b11010111011000;     //118pi/512
   m_cos[118]  =  14'b00110001011100;     //118pi/512
   m_sin[119]  =  14'b11010111000101;     //119pi/512
   m_cos[119]  =  14'b00110001001101;     //119pi/512
   m_sin[120]  =  14'b11010110110011;     //120pi/512
   m_cos[120]  =  14'b00110000111110;     //120pi/512
   m_sin[121]  =  14'b11010110100001;     //121pi/512
   m_cos[121]  =  14'b00110000101110;     //121pi/512
   m_sin[122]  =  14'b11010110001111;     //122pi/512
   m_cos[122]  =  14'b00110000011111;     //122pi/512
   m_sin[123]  =  14'b11010101111100;     //123pi/512
   m_cos[123]  =  14'b00110000001111;     //123pi/512
   m_sin[124]  =  14'b11010101101011;     //124pi/512
   m_cos[124]  =  14'b00101111111111;     //124pi/512
   m_sin[125]  =  14'b11010101011001;     //125pi/512
   m_cos[125]  =  14'b00101111101111;     //125pi/512
   m_sin[126]  =  14'b11010101000111;     //126pi/512
   m_cos[126]  =  14'b00101111011111;     //126pi/512
   m_sin[127]  =  14'b11010100110101;     //127pi/512
   m_cos[127]  =  14'b00101111001111;     //127pi/512
   m_sin[128]  =  14'b11010100100100;     //128pi/512
   m_cos[128]  =  14'b00101110111111;     //128pi/512
   m_sin[129]  =  14'b11010100010010;     //129pi/512
   m_cos[129]  =  14'b00101110101111;     //129pi/512
   m_sin[130]  =  14'b11010100000001;     //130pi/512
   m_cos[130]  =  14'b00101110011111;     //130pi/512
   m_sin[131]  =  14'b11010011101111;     //131pi/512
   m_cos[131]  =  14'b00101110001110;     //131pi/512
   m_sin[132]  =  14'b11010011011110;     //132pi/512
   m_cos[132]  =  14'b00101101111110;     //132pi/512
   m_sin[133]  =  14'b11010011001101;     //133pi/512
   m_cos[133]  =  14'b00101101101101;     //133pi/512
   m_sin[134]  =  14'b11010010111100;     //134pi/512
   m_cos[134]  =  14'b00101101011100;     //134pi/512
   m_sin[135]  =  14'b11010010101011;     //135pi/512
   m_cos[135]  =  14'b00101101001011;     //135pi/512
   m_sin[136]  =  14'b11010010011010;     //136pi/512
   m_cos[136]  =  14'b00101100111010;     //136pi/512
   m_sin[137]  =  14'b11010010001010;     //137pi/512
   m_cos[137]  =  14'b00101100101001;     //137pi/512
   m_sin[138]  =  14'b11010001111001;     //138pi/512
   m_cos[138]  =  14'b00101100011000;     //138pi/512
   m_sin[139]  =  14'b11010001101001;     //139pi/512
   m_cos[139]  =  14'b00101100000111;     //139pi/512
   m_sin[140]  =  14'b11010001011000;     //140pi/512
   m_cos[140]  =  14'b00101011110110;     //140pi/512
   m_sin[141]  =  14'b11010001001000;     //141pi/512
   m_cos[141]  =  14'b00101011100100;     //141pi/512
   m_sin[142]  =  14'b11010000111000;     //142pi/512
   m_cos[142]  =  14'b00101011010011;     //142pi/512
   m_sin[143]  =  14'b11010000101000;     //143pi/512
   m_cos[143]  =  14'b00101011000001;     //143pi/512
   m_sin[144]  =  14'b11010000011000;     //144pi/512
   m_cos[144]  =  14'b00101010101111;     //144pi/512
   m_sin[145]  =  14'b11010000001000;     //145pi/512
   m_cos[145]  =  14'b00101010011101;     //145pi/512
   m_sin[146]  =  14'b11001111111000;     //146pi/512
   m_cos[146]  =  14'b00101010001100;     //146pi/512
   m_sin[147]  =  14'b11001111101000;     //147pi/512
   m_cos[147]  =  14'b00101001111010;     //147pi/512
   m_sin[148]  =  14'b11001111011001;     //148pi/512
   m_cos[148]  =  14'b00101001100111;     //148pi/512
   m_sin[149]  =  14'b11001111001001;     //149pi/512
   m_cos[149]  =  14'b00101001010101;     //149pi/512
   m_sin[150]  =  14'b11001110111010;     //150pi/512
   m_cos[150]  =  14'b00101001000011;     //150pi/512
   m_sin[151]  =  14'b11001110101011;     //151pi/512
   m_cos[151]  =  14'b00101000110001;     //151pi/512
   m_sin[152]  =  14'b11001110011011;     //152pi/512
   m_cos[152]  =  14'b00101000011110;     //152pi/512
   m_sin[153]  =  14'b11001110001100;     //153pi/512
   m_cos[153]  =  14'b00101000001100;     //153pi/512
   m_sin[154]  =  14'b11001101111101;     //154pi/512
   m_cos[154]  =  14'b00100111111001;     //154pi/512
   m_sin[155]  =  14'b11001101101111;     //155pi/512
   m_cos[155]  =  14'b00100111100110;     //155pi/512
   m_sin[156]  =  14'b11001101100000;     //156pi/512
   m_cos[156]  =  14'b00100111010100;     //156pi/512
   m_sin[157]  =  14'b11001101010001;     //157pi/512
   m_cos[157]  =  14'b00100111000001;     //157pi/512
   m_sin[158]  =  14'b11001101000011;     //158pi/512
   m_cos[158]  =  14'b00100110101110;     //158pi/512
   m_sin[159]  =  14'b11001100110100;     //159pi/512
   m_cos[159]  =  14'b00100110011011;     //159pi/512
   m_sin[160]  =  14'b11001100100110;     //160pi/512
   m_cos[160]  =  14'b00100110000111;     //160pi/512
   m_sin[161]  =  14'b11001100011000;     //161pi/512
   m_cos[161]  =  14'b00100101110100;     //161pi/512
   m_sin[162]  =  14'b11001100001010;     //162pi/512
   m_cos[162]  =  14'b00100101100001;     //162pi/512
   m_sin[163]  =  14'b11001011111100;     //163pi/512
   m_cos[163]  =  14'b00100101001110;     //163pi/512
   m_sin[164]  =  14'b11001011101110;     //164pi/512
   m_cos[164]  =  14'b00100100111010;     //164pi/512
   m_sin[165]  =  14'b11001011100000;     //165pi/512
   m_cos[165]  =  14'b00100100100111;     //165pi/512
   m_sin[166]  =  14'b11001011010011;     //166pi/512
   m_cos[166]  =  14'b00100100010011;     //166pi/512
   m_sin[167]  =  14'b11001011000101;     //167pi/512
   m_cos[167]  =  14'b00100011111111;     //167pi/512
   m_sin[168]  =  14'b11001010111000;     //168pi/512
   m_cos[168]  =  14'b00100011101011;     //168pi/512
   m_sin[169]  =  14'b11001010101011;     //169pi/512
   m_cos[169]  =  14'b00100011011000;     //169pi/512
   m_sin[170]  =  14'b11001010011110;     //170pi/512
   m_cos[170]  =  14'b00100011000100;     //170pi/512
   m_sin[171]  =  14'b11001010010000;     //171pi/512
   m_cos[171]  =  14'b00100010110000;     //171pi/512
   m_sin[172]  =  14'b11001010000100;     //172pi/512
   m_cos[172]  =  14'b00100010011100;     //172pi/512
   m_sin[173]  =  14'b11001001110111;     //173pi/512
   m_cos[173]  =  14'b00100010000111;     //173pi/512
   m_sin[174]  =  14'b11001001101010;     //174pi/512
   m_cos[174]  =  14'b00100001110011;     //174pi/512
   m_sin[175]  =  14'b11001001011110;     //175pi/512
   m_cos[175]  =  14'b00100001011111;     //175pi/512
   m_sin[176]  =  14'b11001001010001;     //176pi/512
   m_cos[176]  =  14'b00100001001010;     //176pi/512
   m_sin[177]  =  14'b11001001000101;     //177pi/512
   m_cos[177]  =  14'b00100000110110;     //177pi/512
   m_sin[178]  =  14'b11001000111001;     //178pi/512
   m_cos[178]  =  14'b00100000100010;     //178pi/512
   m_sin[179]  =  14'b11001000101101;     //179pi/512
   m_cos[179]  =  14'b00100000001101;     //179pi/512
   m_sin[180]  =  14'b11001000100001;     //180pi/512
   m_cos[180]  =  14'b00011111111000;     //180pi/512
   m_sin[181]  =  14'b11001000010101;     //181pi/512
   m_cos[181]  =  14'b00011111100100;     //181pi/512
   m_sin[182]  =  14'b11001000001001;     //182pi/512
   m_cos[182]  =  14'b00011111001111;     //182pi/512
   m_sin[183]  =  14'b11000111111101;     //183pi/512
   m_cos[183]  =  14'b00011110111010;     //183pi/512
   m_sin[184]  =  14'b11000111110010;     //184pi/512
   m_cos[184]  =  14'b00011110100101;     //184pi/512
   m_sin[185]  =  14'b11000111100111;     //185pi/512
   m_cos[185]  =  14'b00011110010000;     //185pi/512
   m_sin[186]  =  14'b11000111011011;     //186pi/512
   m_cos[186]  =  14'b00011101111011;     //186pi/512
   m_sin[187]  =  14'b11000111010000;     //187pi/512
   m_cos[187]  =  14'b00011101100110;     //187pi/512
   m_sin[188]  =  14'b11000111000101;     //188pi/512
   m_cos[188]  =  14'b00011101010000;     //188pi/512
   m_sin[189]  =  14'b11000110111010;     //189pi/512
   m_cos[189]  =  14'b00011100111011;     //189pi/512
   m_sin[190]  =  14'b11000110110000;     //190pi/512
   m_cos[190]  =  14'b00011100100110;     //190pi/512
   m_sin[191]  =  14'b11000110100101;     //191pi/512
   m_cos[191]  =  14'b00011100010000;     //191pi/512
   m_sin[192]  =  14'b11000110011011;     //192pi/512
   m_cos[192]  =  14'b00011011111011;     //192pi/512
   m_sin[193]  =  14'b11000110010000;     //193pi/512
   m_cos[193]  =  14'b00011011100110;     //193pi/512
   m_sin[194]  =  14'b11000110000110;     //194pi/512
   m_cos[194]  =  14'b00011011010000;     //194pi/512
   m_sin[195]  =  14'b11000101111100;     //195pi/512
   m_cos[195]  =  14'b00011010111010;     //195pi/512
   m_sin[196]  =  14'b11000101110010;     //196pi/512
   m_cos[196]  =  14'b00011010100101;     //196pi/512
   m_sin[197]  =  14'b11000101101000;     //197pi/512
   m_cos[197]  =  14'b00011010001111;     //197pi/512
   m_sin[198]  =  14'b11000101011110;     //198pi/512
   m_cos[198]  =  14'b00011001111001;     //198pi/512
   m_sin[199]  =  14'b11000101010101;     //199pi/512
   m_cos[199]  =  14'b00011001100011;     //199pi/512
   m_sin[200]  =  14'b11000101001011;     //200pi/512
   m_cos[200]  =  14'b00011001001101;     //200pi/512
   m_sin[201]  =  14'b11000101000010;     //201pi/512
   m_cos[201]  =  14'b00011000110111;     //201pi/512
   m_sin[202]  =  14'b11000100111001;     //202pi/512
   m_cos[202]  =  14'b00011000100001;     //202pi/512
   m_sin[203]  =  14'b11000100110000;     //203pi/512
   m_cos[203]  =  14'b00011000001011;     //203pi/512
   m_sin[204]  =  14'b11000100100111;     //204pi/512
   m_cos[204]  =  14'b00010111110101;     //204pi/512
   m_sin[205]  =  14'b11000100011110;     //205pi/512
   m_cos[205]  =  14'b00010111011111;     //205pi/512
   m_sin[206]  =  14'b11000100010101;     //206pi/512
   m_cos[206]  =  14'b00010111001001;     //206pi/512
   m_sin[207]  =  14'b11000100001101;     //207pi/512
   m_cos[207]  =  14'b00010110110010;     //207pi/512
   m_sin[208]  =  14'b11000100000100;     //208pi/512
   m_cos[208]  =  14'b00010110011100;     //208pi/512
   m_sin[209]  =  14'b11000011111100;     //209pi/512
   m_cos[209]  =  14'b00010110000110;     //209pi/512
   m_sin[210]  =  14'b11000011110100;     //210pi/512
   m_cos[210]  =  14'b00010101101111;     //210pi/512
   m_sin[211]  =  14'b11000011101100;     //211pi/512
   m_cos[211]  =  14'b00010101011001;     //211pi/512
   m_sin[212]  =  14'b11000011100100;     //212pi/512
   m_cos[212]  =  14'b00010101000010;     //212pi/512
   m_sin[213]  =  14'b11000011011100;     //213pi/512
   m_cos[213]  =  14'b00010100101100;     //213pi/512
   m_sin[214]  =  14'b11000011010100;     //214pi/512
   m_cos[214]  =  14'b00010100010101;     //214pi/512
   m_sin[215]  =  14'b11000011001101;     //215pi/512
   m_cos[215]  =  14'b00010011111110;     //215pi/512
   m_sin[216]  =  14'b11000011000101;     //216pi/512
   m_cos[216]  =  14'b00010011101000;     //216pi/512
   m_sin[217]  =  14'b11000010111110;     //217pi/512
   m_cos[217]  =  14'b00010011010001;     //217pi/512
   m_sin[218]  =  14'b11000010110111;     //218pi/512
   m_cos[218]  =  14'b00010010111010;     //218pi/512
   m_sin[219]  =  14'b11000010110000;     //219pi/512
   m_cos[219]  =  14'b00010010100011;     //219pi/512
   m_sin[220]  =  14'b11000010101001;     //220pi/512
   m_cos[220]  =  14'b00010010001100;     //220pi/512
   m_sin[221]  =  14'b11000010100010;     //221pi/512
   m_cos[221]  =  14'b00010001110110;     //221pi/512
   m_sin[222]  =  14'b11000010011100;     //222pi/512
   m_cos[222]  =  14'b00010001011111;     //222pi/512
   m_sin[223]  =  14'b11000010010101;     //223pi/512
   m_cos[223]  =  14'b00010001001000;     //223pi/512
   m_sin[224]  =  14'b11000010001111;     //224pi/512
   m_cos[224]  =  14'b00010000110001;     //224pi/512
   m_sin[225]  =  14'b11000010001001;     //225pi/512
   m_cos[225]  =  14'b00010000011010;     //225pi/512
   m_sin[226]  =  14'b11000010000011;     //226pi/512
   m_cos[226]  =  14'b00010000000010;     //226pi/512
   m_sin[227]  =  14'b11000001111101;     //227pi/512
   m_cos[227]  =  14'b00001111101011;     //227pi/512
   m_sin[228]  =  14'b11000001110111;     //228pi/512
   m_cos[228]  =  14'b00001111010100;     //228pi/512
   m_sin[229]  =  14'b11000001110001;     //229pi/512
   m_cos[229]  =  14'b00001110111101;     //229pi/512
   m_sin[230]  =  14'b11000001101100;     //230pi/512
   m_cos[230]  =  14'b00001110100110;     //230pi/512
   m_sin[231]  =  14'b11000001100111;     //231pi/512
   m_cos[231]  =  14'b00001110001110;     //231pi/512
   m_sin[232]  =  14'b11000001100001;     //232pi/512
   m_cos[232]  =  14'b00001101110111;     //232pi/512
   m_sin[233]  =  14'b11000001011100;     //233pi/512
   m_cos[233]  =  14'b00001101100000;     //233pi/512
   m_sin[234]  =  14'b11000001010111;     //234pi/512
   m_cos[234]  =  14'b00001101001000;     //234pi/512
   m_sin[235]  =  14'b11000001010010;     //235pi/512
   m_cos[235]  =  14'b00001100110001;     //235pi/512
   m_sin[236]  =  14'b11000001001110;     //236pi/512
   m_cos[236]  =  14'b00001100011010;     //236pi/512
   m_sin[237]  =  14'b11000001001001;     //237pi/512
   m_cos[237]  =  14'b00001100000010;     //237pi/512
   m_sin[238]  =  14'b11000001000101;     //238pi/512
   m_cos[238]  =  14'b00001011101011;     //238pi/512
   m_sin[239]  =  14'b11000001000000;     //239pi/512
   m_cos[239]  =  14'b00001011010011;     //239pi/512
   m_sin[240]  =  14'b11000000111100;     //240pi/512
   m_cos[240]  =  14'b00001010111100;     //240pi/512
   m_sin[241]  =  14'b11000000111000;     //241pi/512
   m_cos[241]  =  14'b00001010100100;     //241pi/512
   m_sin[242]  =  14'b11000000110100;     //242pi/512
   m_cos[242]  =  14'b00001010001101;     //242pi/512
   m_sin[243]  =  14'b11000000110001;     //243pi/512
   m_cos[243]  =  14'b00001001110101;     //243pi/512
   m_sin[244]  =  14'b11000000101101;     //244pi/512
   m_cos[244]  =  14'b00001001011101;     //244pi/512
   m_sin[245]  =  14'b11000000101010;     //245pi/512
   m_cos[245]  =  14'b00001001000110;     //245pi/512
   m_sin[246]  =  14'b11000000100110;     //246pi/512
   m_cos[246]  =  14'b00001000101110;     //246pi/512
   m_sin[247]  =  14'b11000000100011;     //247pi/512
   m_cos[247]  =  14'b00001000010111;     //247pi/512
   m_sin[248]  =  14'b11000000100000;     //248pi/512
   m_cos[248]  =  14'b00000111111111;     //248pi/512
   m_sin[249]  =  14'b11000000011101;     //249pi/512
   m_cos[249]  =  14'b00000111100111;     //249pi/512
   m_sin[250]  =  14'b11000000011010;     //250pi/512
   m_cos[250]  =  14'b00000111001111;     //250pi/512
   m_sin[251]  =  14'b11000000011000;     //251pi/512
   m_cos[251]  =  14'b00000110111000;     //251pi/512
   m_sin[252]  =  14'b11000000010101;     //252pi/512
   m_cos[252]  =  14'b00000110100000;     //252pi/512
   m_sin[253]  =  14'b11000000010011;     //253pi/512
   m_cos[253]  =  14'b00000110001000;     //253pi/512
   m_sin[254]  =  14'b11000000010001;     //254pi/512
   m_cos[254]  =  14'b00000101110000;     //254pi/512
   m_sin[255]  =  14'b11000000001111;     //255pi/512
   m_cos[255]  =  14'b00000101011001;     //255pi/512
   m_sin[256]  =  14'b11000000001101;     //256pi/512
   m_cos[256]  =  14'b00000101000001;     //256pi/512
   m_sin[257]  =  14'b11000000001011;     //257pi/512
   m_cos[257]  =  14'b00000100101001;     //257pi/512
   m_sin[258]  =  14'b11000000001001;     //258pi/512
   m_cos[258]  =  14'b00000100010001;     //258pi/512
   m_sin[259]  =  14'b11000000001000;     //259pi/512
   m_cos[259]  =  14'b00000011111001;     //259pi/512
   m_sin[260]  =  14'b11000000000110;     //260pi/512
   m_cos[260]  =  14'b00000011100010;     //260pi/512
   m_sin[261]  =  14'b11000000000101;     //261pi/512
   m_cos[261]  =  14'b00000011001010;     //261pi/512
   m_sin[262]  =  14'b11000000000100;     //262pi/512
   m_cos[262]  =  14'b00000010110010;     //262pi/512
   m_sin[263]  =  14'b11000000000011;     //263pi/512
   m_cos[263]  =  14'b00000010011010;     //263pi/512
   m_sin[264]  =  14'b11000000000010;     //264pi/512
   m_cos[264]  =  14'b00000010000010;     //264pi/512
   m_sin[265]  =  14'b11000000000001;     //265pi/512
   m_cos[265]  =  14'b00000001101010;     //265pi/512
   m_sin[266]  =  14'b11000000000001;     //266pi/512
   m_cos[266]  =  14'b00000001010010;     //266pi/512
   m_sin[267]  =  14'b11000000000000;     //267pi/512
   m_cos[267]  =  14'b00000000111011;     //267pi/512
   m_sin[268]  =  14'b11000000000000;     //268pi/512
   m_cos[268]  =  14'b00000000100011;     //268pi/512
   m_sin[269]  =  14'b11000000000000;     //269pi/512
   m_cos[269]  =  14'b00000000001011;     //269pi/512
   m_sin[270]  =  14'b11000000000000;     //270pi/512
   m_cos[270]  =  14'b11111111110011;     //270pi/512
   m_sin[271]  =  14'b11000000000000;     //271pi/512
   m_cos[271]  =  14'b11111111011100;     //271pi/512
   m_sin[272]  =  14'b11000000000000;     //272pi/512
   m_cos[272]  =  14'b11111111000100;     //272pi/512
   m_sin[273]  =  14'b11000000000001;     //273pi/512
   m_cos[273]  =  14'b11111110101100;     //273pi/512
   m_sin[274]  =  14'b11000000000001;     //274pi/512
   m_cos[274]  =  14'b11111110010100;     //274pi/512
   m_sin[275]  =  14'b11000000000010;     //275pi/512
   m_cos[275]  =  14'b11111101111100;     //275pi/512
   m_sin[276]  =  14'b11000000000011;     //276pi/512
   m_cos[276]  =  14'b11111101100100;     //276pi/512
   m_sin[277]  =  14'b11000000000100;     //277pi/512
   m_cos[277]  =  14'b11111101001100;     //277pi/512
   m_sin[278]  =  14'b11000000000101;     //278pi/512
   m_cos[278]  =  14'b11111100110101;     //278pi/512
   m_sin[279]  =  14'b11000000000110;     //279pi/512
   m_cos[279]  =  14'b11111100011101;     //279pi/512
   m_sin[280]  =  14'b11000000001000;     //280pi/512
   m_cos[280]  =  14'b11111100000101;     //280pi/512
   m_sin[281]  =  14'b11000000001001;     //281pi/512
   m_cos[281]  =  14'b11111011101101;     //281pi/512
   m_sin[282]  =  14'b11000000001011;     //282pi/512
   m_cos[282]  =  14'b11111011010101;     //282pi/512
   m_sin[283]  =  14'b11000000001101;     //283pi/512
   m_cos[283]  =  14'b11111010111101;     //283pi/512
   m_sin[284]  =  14'b11000000001111;     //284pi/512
   m_cos[284]  =  14'b11111010100110;     //284pi/512
   m_sin[285]  =  14'b11000000010001;     //285pi/512
   m_cos[285]  =  14'b11111010001110;     //285pi/512
   m_sin[286]  =  14'b11000000010011;     //286pi/512
   m_cos[286]  =  14'b11111001110110;     //286pi/512
   m_sin[287]  =  14'b11000000010101;     //287pi/512
   m_cos[287]  =  14'b11111001011110;     //287pi/512
   m_sin[288]  =  14'b11000000011000;     //288pi/512
   m_cos[288]  =  14'b11111001000111;     //288pi/512
   m_sin[289]  =  14'b11000000011011;     //289pi/512
   m_cos[289]  =  14'b11111000101111;     //289pi/512
   m_sin[290]  =  14'b11000000011101;     //290pi/512
   m_cos[290]  =  14'b11111000010111;     //290pi/512
   m_sin[291]  =  14'b11000000100000;     //291pi/512
   m_cos[291]  =  14'b11110111111111;     //291pi/512
   m_sin[292]  =  14'b11000000100011;     //292pi/512
   m_cos[292]  =  14'b11110111101000;     //292pi/512
   m_sin[293]  =  14'b11000000100110;     //293pi/512
   m_cos[293]  =  14'b11110111010000;     //293pi/512
   m_sin[294]  =  14'b11000000101010;     //294pi/512
   m_cos[294]  =  14'b11110110111000;     //294pi/512
   m_sin[295]  =  14'b11000000101101;     //295pi/512
   m_cos[295]  =  14'b11110110100001;     //295pi/512
   m_sin[296]  =  14'b11000000110001;     //296pi/512
   m_cos[296]  =  14'b11110110001001;     //296pi/512
   m_sin[297]  =  14'b11000000110101;     //297pi/512
   m_cos[297]  =  14'b11110101110010;     //297pi/512
   m_sin[298]  =  14'b11000000111000;     //298pi/512
   m_cos[298]  =  14'b11110101011010;     //298pi/512
   m_sin[299]  =  14'b11000000111101;     //299pi/512
   m_cos[299]  =  14'b11110101000011;     //299pi/512
   m_sin[300]  =  14'b11000001000001;     //300pi/512
   m_cos[300]  =  14'b11110100101011;     //300pi/512
   m_sin[301]  =  14'b11000001000101;     //301pi/512
   m_cos[301]  =  14'b11110100010100;     //301pi/512
   m_sin[302]  =  14'b11000001001001;     //302pi/512
   m_cos[302]  =  14'b11110011111100;     //302pi/512
   m_sin[303]  =  14'b11000001001110;     //303pi/512
   m_cos[303]  =  14'b11110011100101;     //303pi/512
   m_sin[304]  =  14'b11000001010011;     //304pi/512
   m_cos[304]  =  14'b11110011001101;     //304pi/512
   m_sin[305]  =  14'b11000001011000;     //305pi/512
   m_cos[305]  =  14'b11110010110110;     //305pi/512
   m_sin[306]  =  14'b11000001011100;     //306pi/512
   m_cos[306]  =  14'b11110010011110;     //306pi/512
   m_sin[307]  =  14'b11000001100010;     //307pi/512
   m_cos[307]  =  14'b11110010000111;     //307pi/512
   m_sin[308]  =  14'b11000001100111;     //308pi/512
   m_cos[308]  =  14'b11110001110000;     //308pi/512
   m_sin[309]  =  14'b11000001101100;     //309pi/512
   m_cos[309]  =  14'b11110001011001;     //309pi/512
   m_sin[310]  =  14'b11000001110010;     //310pi/512
   m_cos[310]  =  14'b11110001000001;     //310pi/512
   m_sin[311]  =  14'b11000001110111;     //311pi/512
   m_cos[311]  =  14'b11110000101010;     //311pi/512
   m_sin[312]  =  14'b11000001111101;     //312pi/512
   m_cos[312]  =  14'b11110000010011;     //312pi/512
   m_sin[313]  =  14'b11000010000011;     //313pi/512
   m_cos[313]  =  14'b11101111111100;     //313pi/512
   m_sin[314]  =  14'b11000010001001;     //314pi/512
   m_cos[314]  =  14'b11101111100101;     //314pi/512
   m_sin[315]  =  14'b11000010001111;     //315pi/512
   m_cos[315]  =  14'b11101111001110;     //315pi/512
   m_sin[316]  =  14'b11000010010110;     //316pi/512
   m_cos[316]  =  14'b11101110110111;     //316pi/512
   m_sin[317]  =  14'b11000010011100;     //317pi/512
   m_cos[317]  =  14'b11101110100000;     //317pi/512
   m_sin[318]  =  14'b11000010100011;     //318pi/512
   m_cos[318]  =  14'b11101110001001;     //318pi/512
   m_sin[319]  =  14'b11000010101010;     //319pi/512
   m_cos[319]  =  14'b11101101110010;     //319pi/512
   m_sin[320]  =  14'b11000010110000;     //320pi/512
   m_cos[320]  =  14'b11101101011011;     //320pi/512
   m_sin[321]  =  14'b11000010110111;     //321pi/512
   m_cos[321]  =  14'b11101101000100;     //321pi/512
   m_sin[322]  =  14'b11000010111111;     //322pi/512
   m_cos[322]  =  14'b11101100101101;     //322pi/512
   m_sin[323]  =  14'b11000011000110;     //323pi/512
   m_cos[323]  =  14'b11101100010111;     //323pi/512
   m_sin[324]  =  14'b11000011001101;     //324pi/512
   m_cos[324]  =  14'b11101100000000;     //324pi/512
   m_sin[325]  =  14'b11000011010101;     //325pi/512
   m_cos[325]  =  14'b11101011101001;     //325pi/512
   m_sin[326]  =  14'b11000011011100;     //326pi/512
   m_cos[326]  =  14'b11101011010011;     //326pi/512
   m_sin[327]  =  14'b11000011100100;     //327pi/512
   m_cos[327]  =  14'b11101010111100;     //327pi/512
   m_sin[328]  =  14'b11000011101100;     //328pi/512
   m_cos[328]  =  14'b11101010100110;     //328pi/512
   m_sin[329]  =  14'b11000011110100;     //329pi/512
   m_cos[329]  =  14'b11101010001111;     //329pi/512
   m_sin[330]  =  14'b11000011111100;     //330pi/512
   m_cos[330]  =  14'b11101001111001;     //330pi/512
   m_sin[331]  =  14'b11000100000101;     //331pi/512
   m_cos[331]  =  14'b11101001100010;     //331pi/512
   m_sin[332]  =  14'b11000100001101;     //332pi/512
   m_cos[332]  =  14'b11101001001100;     //332pi/512
   m_sin[333]  =  14'b11000100010110;     //333pi/512
   m_cos[333]  =  14'b11101000110110;     //333pi/512
   m_sin[334]  =  14'b11000100011110;     //334pi/512
   m_cos[334]  =  14'b11101000011111;     //334pi/512
   m_sin[335]  =  14'b11000100100111;     //335pi/512
   m_cos[335]  =  14'b11101000001001;     //335pi/512
   m_sin[336]  =  14'b11000100110000;     //336pi/512
   m_cos[336]  =  14'b11100111110011;     //336pi/512
   m_sin[337]  =  14'b11000100111001;     //337pi/512
   m_cos[337]  =  14'b11100111011101;     //337pi/512
   m_sin[338]  =  14'b11000101000010;     //338pi/512
   m_cos[338]  =  14'b11100111000111;     //338pi/512
   m_sin[339]  =  14'b11000101001100;     //339pi/512
   m_cos[339]  =  14'b11100110110001;     //339pi/512
   m_sin[340]  =  14'b11000101010101;     //340pi/512
   m_cos[340]  =  14'b11100110011011;     //340pi/512
   m_sin[341]  =  14'b11000101011111;     //341pi/512
   m_cos[341]  =  14'b11100110000101;     //341pi/512
   m_sin[342]  =  14'b11000101101001;     //342pi/512
   m_cos[342]  =  14'b11100101101111;     //342pi/512
   m_sin[343]  =  14'b11000101110010;     //343pi/512
   m_cos[343]  =  14'b11100101011010;     //343pi/512
   m_sin[344]  =  14'b11000101111100;     //344pi/512
   m_cos[344]  =  14'b11100101000100;     //344pi/512
   m_sin[345]  =  14'b11000110000111;     //345pi/512
   m_cos[345]  =  14'b11100100101110;     //345pi/512
   m_sin[346]  =  14'b11000110010001;     //346pi/512
   m_cos[346]  =  14'b11100100011001;     //346pi/512
   m_sin[347]  =  14'b11000110011011;     //347pi/512
   m_cos[347]  =  14'b11100100000011;     //347pi/512
   m_sin[348]  =  14'b11000110100110;     //348pi/512
   m_cos[348]  =  14'b11100011101110;     //348pi/512
   m_sin[349]  =  14'b11000110110000;     //349pi/512
   m_cos[349]  =  14'b11100011011001;     //349pi/512
   m_sin[350]  =  14'b11000110111011;     //350pi/512
   m_cos[350]  =  14'b11100011000011;     //350pi/512
   m_sin[351]  =  14'b11000111000110;     //351pi/512
   m_cos[351]  =  14'b11100010101110;     //351pi/512
   m_sin[352]  =  14'b11000111010001;     //352pi/512
   m_cos[352]  =  14'b11100010011001;     //352pi/512
   m_sin[353]  =  14'b11000111011100;     //353pi/512
   m_cos[353]  =  14'b11100010000100;     //353pi/512
   m_sin[354]  =  14'b11000111100111;     //354pi/512
   m_cos[354]  =  14'b11100001101111;     //354pi/512
   m_sin[355]  =  14'b11000111110011;     //355pi/512
   m_cos[355]  =  14'b11100001011010;     //355pi/512
   m_sin[356]  =  14'b11000111111110;     //356pi/512
   m_cos[356]  =  14'b11100001000101;     //356pi/512
   m_sin[357]  =  14'b11001000001010;     //357pi/512
   m_cos[357]  =  14'b11100000110000;     //357pi/512
   m_sin[358]  =  14'b11001000010101;     //358pi/512
   m_cos[358]  =  14'b11100000011011;     //358pi/512
   m_sin[359]  =  14'b11001000100001;     //359pi/512
   m_cos[359]  =  14'b11100000000110;     //359pi/512
   m_sin[360]  =  14'b11001000101101;     //360pi/512
   m_cos[360]  =  14'b11011111110010;     //360pi/512
   m_sin[361]  =  14'b11001000111001;     //361pi/512
   m_cos[361]  =  14'b11011111011101;     //361pi/512
   m_sin[362]  =  14'b11001001000101;     //362pi/512
   m_cos[362]  =  14'b11011111001000;     //362pi/512
   m_sin[363]  =  14'b11001001010010;     //363pi/512
   m_cos[363]  =  14'b11011110110100;     //363pi/512
   m_sin[364]  =  14'b11001001011110;     //364pi/512
   m_cos[364]  =  14'b11011110100000;     //364pi/512
   m_sin[365]  =  14'b11001001101011;     //365pi/512
   m_cos[365]  =  14'b11011110001011;     //365pi/512
   m_sin[366]  =  14'b11001001110111;     //366pi/512
   m_cos[366]  =  14'b11011101110111;     //366pi/512
   m_sin[367]  =  14'b11001010000100;     //367pi/512
   m_cos[367]  =  14'b11011101100011;     //367pi/512
   m_sin[368]  =  14'b11001010010001;     //368pi/512
   m_cos[368]  =  14'b11011101001111;     //368pi/512
   m_sin[369]  =  14'b11001010011110;     //369pi/512
   m_cos[369]  =  14'b11011100111011;     //369pi/512
   m_sin[370]  =  14'b11001010101011;     //370pi/512
   m_cos[370]  =  14'b11011100100111;     //370pi/512
   m_sin[371]  =  14'b11001010111001;     //371pi/512
   m_cos[371]  =  14'b11011100010011;     //371pi/512
   m_sin[372]  =  14'b11001011000110;     //372pi/512
   m_cos[372]  =  14'b11011011111111;     //372pi/512
   m_sin[373]  =  14'b11001011010011;     //373pi/512
   m_cos[373]  =  14'b11011011101100;     //373pi/512
   m_sin[374]  =  14'b11001011100001;     //374pi/512
   m_cos[374]  =  14'b11011011011000;     //374pi/512
   m_sin[375]  =  14'b11001011101111;     //375pi/512
   m_cos[375]  =  14'b11011011000100;     //375pi/512
   m_sin[376]  =  14'b11001011111101;     //376pi/512
   m_cos[376]  =  14'b11011010110001;     //376pi/512
   m_sin[377]  =  14'b11001100001011;     //377pi/512
   m_cos[377]  =  14'b11011010011110;     //377pi/512
   m_sin[378]  =  14'b11001100011001;     //378pi/512
   m_cos[378]  =  14'b11011010001010;     //378pi/512
   m_sin[379]  =  14'b11001100100111;     //379pi/512
   m_cos[379]  =  14'b11011001110111;     //379pi/512
   m_sin[380]  =  14'b11001100110101;     //380pi/512
   m_cos[380]  =  14'b11011001100100;     //380pi/512
   m_sin[381]  =  14'b11001101000011;     //381pi/512
   m_cos[381]  =  14'b11011001010001;     //381pi/512
   m_sin[382]  =  14'b11001101010010;     //382pi/512
   m_cos[382]  =  14'b11011000111110;     //382pi/512
   m_sin[383]  =  14'b11001101100001;     //383pi/512
   m_cos[383]  =  14'b11011000101011;     //383pi/512
   m_sin[384]  =  14'b11001101101111;     //384pi/512
   m_cos[384]  =  14'b11011000011000;     //384pi/512
   m_sin[385]  =  14'b11001101111110;     //385pi/512
   m_cos[385]  =  14'b11011000000101;     //385pi/512
   m_sin[386]  =  14'b11001110001101;     //386pi/512
   m_cos[386]  =  14'b11010111110011;     //386pi/512
   m_sin[387]  =  14'b11001110011100;     //387pi/512
   m_cos[387]  =  14'b11010111100000;     //387pi/512
   m_sin[388]  =  14'b11001110101011;     //388pi/512
   m_cos[388]  =  14'b11010111001110;     //388pi/512
   m_sin[389]  =  14'b11001110111011;     //389pi/512
   m_cos[389]  =  14'b11010110111100;     //389pi/512
   m_sin[390]  =  14'b11001111001010;     //390pi/512
   m_cos[390]  =  14'b11010110101001;     //390pi/512
   m_sin[391]  =  14'b11001111011001;     //391pi/512
   m_cos[391]  =  14'b11010110010111;     //391pi/512
   m_sin[392]  =  14'b11001111101001;     //392pi/512
   m_cos[392]  =  14'b11010110000101;     //392pi/512
   m_sin[393]  =  14'b11001111111001;     //393pi/512
   m_cos[393]  =  14'b11010101110011;     //393pi/512
   m_sin[394]  =  14'b11010000001001;     //394pi/512
   m_cos[394]  =  14'b11010101100001;     //394pi/512
   m_sin[395]  =  14'b11010000011000;     //395pi/512
   m_cos[395]  =  14'b11010101001111;     //395pi/512
   m_sin[396]  =  14'b11010000101000;     //396pi/512
   m_cos[396]  =  14'b11010100111110;     //396pi/512
   m_sin[397]  =  14'b11010000111001;     //397pi/512
   m_cos[397]  =  14'b11010100101100;     //397pi/512
   m_sin[398]  =  14'b11010001001001;     //398pi/512
   m_cos[398]  =  14'b11010100011010;     //398pi/512
   m_sin[399]  =  14'b11010001011001;     //399pi/512
   m_cos[399]  =  14'b11010100001001;     //399pi/512
   m_sin[400]  =  14'b11010001101001;     //400pi/512
   m_cos[400]  =  14'b11010011111000;     //400pi/512
   m_sin[401]  =  14'b11010001111010;     //401pi/512
   m_cos[401]  =  14'b11010011100110;     //401pi/512
   m_sin[402]  =  14'b11010010001011;     //402pi/512
   m_cos[402]  =  14'b11010011010101;     //402pi/512
   m_sin[403]  =  14'b11010010011011;     //403pi/512
   m_cos[403]  =  14'b11010011000100;     //403pi/512
   m_sin[404]  =  14'b11010010101100;     //404pi/512
   m_cos[404]  =  14'b11010010110011;     //404pi/512
   m_sin[405]  =  14'b11010010111101;     //405pi/512
   m_cos[405]  =  14'b11010010100010;     //405pi/512
   m_sin[406]  =  14'b11010011001110;     //406pi/512
   m_cos[406]  =  14'b11010010010010;     //406pi/512
   m_sin[407]  =  14'b11010011011111;     //407pi/512
   m_cos[407]  =  14'b11010010000001;     //407pi/512
   m_sin[408]  =  14'b11010011110000;     //408pi/512
   m_cos[408]  =  14'b11010001110000;     //408pi/512
   m_sin[409]  =  14'b11010100000010;     //409pi/512
   m_cos[409]  =  14'b11010001100000;     //409pi/512
   m_sin[410]  =  14'b11010100010011;     //410pi/512
   m_cos[410]  =  14'b11010001010000;     //410pi/512
   m_sin[411]  =  14'b11010100100101;     //411pi/512
   m_cos[411]  =  14'b11010000111111;     //411pi/512
   m_sin[412]  =  14'b11010100110110;     //412pi/512
   m_cos[412]  =  14'b11010000101111;     //412pi/512
   m_sin[413]  =  14'b11010101001000;     //413pi/512
   m_cos[413]  =  14'b11010000011111;     //413pi/512
   m_sin[414]  =  14'b11010101011010;     //414pi/512
   m_cos[414]  =  14'b11010000001111;     //414pi/512
   m_sin[415]  =  14'b11010101101011;     //415pi/512
   m_cos[415]  =  14'b11001111111111;     //415pi/512
   m_sin[416]  =  14'b11010101111101;     //416pi/512
   m_cos[416]  =  14'b11001111110000;     //416pi/512
   m_sin[417]  =  14'b11010110001111;     //417pi/512
   m_cos[417]  =  14'b11001111100000;     //417pi/512
   m_sin[418]  =  14'b11010110100010;     //418pi/512
   m_cos[418]  =  14'b11001111010000;     //418pi/512
   m_sin[419]  =  14'b11010110110100;     //419pi/512
   m_cos[419]  =  14'b11001111000001;     //419pi/512
   m_sin[420]  =  14'b11010111000110;     //420pi/512
   m_cos[420]  =  14'b11001110110010;     //420pi/512
   m_sin[421]  =  14'b11010111011001;     //421pi/512
   m_cos[421]  =  14'b11001110100011;     //421pi/512
   m_sin[422]  =  14'b11010111101011;     //422pi/512
   m_cos[422]  =  14'b11001110010011;     //422pi/512
   m_sin[423]  =  14'b11010111111110;     //423pi/512
   m_cos[423]  =  14'b11001110000100;     //423pi/512
   m_sin[424]  =  14'b11011000010000;     //424pi/512
   m_cos[424]  =  14'b11001101110110;     //424pi/512
   m_sin[425]  =  14'b11011000100011;     //425pi/512
   m_cos[425]  =  14'b11001101100111;     //425pi/512
   m_sin[426]  =  14'b11011000110110;     //426pi/512
   m_cos[426]  =  14'b11001101011000;     //426pi/512
   m_sin[427]  =  14'b11011001001001;     //427pi/512
   m_cos[427]  =  14'b11001101001010;     //427pi/512
   m_sin[428]  =  14'b11011001011100;     //428pi/512
   m_cos[428]  =  14'b11001100111011;     //428pi/512
   m_sin[429]  =  14'b11011001101111;     //429pi/512
   m_cos[429]  =  14'b11001100101101;     //429pi/512
   m_sin[430]  =  14'b11011010000010;     //430pi/512
   m_cos[430]  =  14'b11001100011111;     //430pi/512
   m_sin[431]  =  14'b11011010010101;     //431pi/512
   m_cos[431]  =  14'b11001100010000;     //431pi/512
   m_sin[432]  =  14'b11011010101001;     //432pi/512
   m_cos[432]  =  14'b11001100000010;     //432pi/512
   m_sin[433]  =  14'b11011010111100;     //433pi/512
   m_cos[433]  =  14'b11001011110101;     //433pi/512
   m_sin[434]  =  14'b11011011010000;     //434pi/512
   m_cos[434]  =  14'b11001011100111;     //434pi/512
   m_sin[435]  =  14'b11011011100011;     //435pi/512
   m_cos[435]  =  14'b11001011011001;     //435pi/512
   m_sin[436]  =  14'b11011011110111;     //436pi/512
   m_cos[436]  =  14'b11001011001100;     //436pi/512
   m_sin[437]  =  14'b11011100001011;     //437pi/512
   m_cos[437]  =  14'b11001010111110;     //437pi/512
   m_sin[438]  =  14'b11011100011110;     //438pi/512
   m_cos[438]  =  14'b11001010110001;     //438pi/512
   m_sin[439]  =  14'b11011100110010;     //439pi/512
   m_cos[439]  =  14'b11001010100100;     //439pi/512
   m_sin[440]  =  14'b11011101000110;     //440pi/512
   m_cos[440]  =  14'b11001010010111;     //440pi/512
   m_sin[441]  =  14'b11011101011010;     //441pi/512
   m_cos[441]  =  14'b11001010001010;     //441pi/512
   m_sin[442]  =  14'b11011101101111;     //442pi/512
   m_cos[442]  =  14'b11001001111101;     //442pi/512
   m_sin[443]  =  14'b11011110000011;     //443pi/512
   m_cos[443]  =  14'b11001001110000;     //443pi/512
   m_sin[444]  =  14'b11011110010111;     //444pi/512
   m_cos[444]  =  14'b11001001100011;     //444pi/512
   m_sin[445]  =  14'b11011110101011;     //445pi/512
   m_cos[445]  =  14'b11001001010111;     //445pi/512
   m_sin[446]  =  14'b11011111000000;     //446pi/512
   m_cos[446]  =  14'b11001001001011;     //446pi/512
   m_sin[447]  =  14'b11011111010100;     //447pi/512
   m_cos[447]  =  14'b11001000111110;     //447pi/512
   m_sin[448]  =  14'b11011111101001;     //448pi/512
   m_cos[448]  =  14'b11001000110010;     //448pi/512
   m_sin[449]  =  14'b11011111111101;     //449pi/512
   m_cos[449]  =  14'b11001000100110;     //449pi/512
   m_sin[450]  =  14'b11100000010010;     //450pi/512
   m_cos[450]  =  14'b11001000011010;     //450pi/512
   m_sin[451]  =  14'b11100000100111;     //451pi/512
   m_cos[451]  =  14'b11001000001111;     //451pi/512
   m_sin[452]  =  14'b11100000111100;     //452pi/512
   m_cos[452]  =  14'b11001000000011;     //452pi/512
   m_sin[453]  =  14'b11100001010001;     //453pi/512
   m_cos[453]  =  14'b11000111110111;     //453pi/512
   m_sin[454]  =  14'b11100001100110;     //454pi/512
   m_cos[454]  =  14'b11000111101100;     //454pi/512
   m_sin[455]  =  14'b11100001111011;     //455pi/512
   m_cos[455]  =  14'b11000111100001;     //455pi/512
   m_sin[456]  =  14'b11100010010000;     //456pi/512
   m_cos[456]  =  14'b11000111010110;     //456pi/512
   m_sin[457]  =  14'b11100010100101;     //457pi/512
   m_cos[457]  =  14'b11000111001010;     //457pi/512
   m_sin[458]  =  14'b11100010111010;     //458pi/512
   m_cos[458]  =  14'b11000111000000;     //458pi/512
   m_sin[459]  =  14'b11100011010000;     //459pi/512
   m_cos[459]  =  14'b11000110110101;     //459pi/512
   m_sin[460]  =  14'b11100011100101;     //460pi/512
   m_cos[460]  =  14'b11000110101010;     //460pi/512
   m_sin[461]  =  14'b11100011111010;     //461pi/512
   m_cos[461]  =  14'b11000110100000;     //461pi/512
   m_sin[462]  =  14'b11100100010000;     //462pi/512
   m_cos[462]  =  14'b11000110010101;     //462pi/512
   m_sin[463]  =  14'b11100100100101;     //463pi/512
   m_cos[463]  =  14'b11000110001011;     //463pi/512
   m_sin[464]  =  14'b11100100111011;     //464pi/512
   m_cos[464]  =  14'b11000110000001;     //464pi/512
   m_sin[465]  =  14'b11100101010001;     //465pi/512
   m_cos[465]  =  14'b11000101110111;     //465pi/512
   m_sin[466]  =  14'b11100101100110;     //466pi/512
   m_cos[466]  =  14'b11000101101101;     //466pi/512
   m_sin[467]  =  14'b11100101111100;     //467pi/512
   m_cos[467]  =  14'b11000101100011;     //467pi/512
   m_sin[468]  =  14'b11100110010010;     //468pi/512
   m_cos[468]  =  14'b11000101011001;     //468pi/512
   m_sin[469]  =  14'b11100110101000;     //469pi/512
   m_cos[469]  =  14'b11000101010000;     //469pi/512
   m_sin[470]  =  14'b11100110111110;     //470pi/512
   m_cos[470]  =  14'b11000101000110;     //470pi/512
   m_sin[471]  =  14'b11100111010100;     //471pi/512
   m_cos[471]  =  14'b11000100111101;     //471pi/512
   m_sin[472]  =  14'b11100111101010;     //472pi/512
   m_cos[472]  =  14'b11000100110100;     //472pi/512
   m_sin[473]  =  14'b11101000000000;     //473pi/512
   m_cos[473]  =  14'b11000100101011;     //473pi/512
   m_sin[474]  =  14'b11101000010110;     //474pi/512
   m_cos[474]  =  14'b11000100100010;     //474pi/512
   m_sin[475]  =  14'b11101000101100;     //475pi/512
   m_cos[475]  =  14'b11000100011001;     //475pi/512
   m_sin[476]  =  14'b11101001000011;     //476pi/512
   m_cos[476]  =  14'b11000100010001;     //476pi/512
   m_sin[477]  =  14'b11101001011001;     //477pi/512
   m_cos[477]  =  14'b11000100001000;     //477pi/512
   m_sin[478]  =  14'b11101001101111;     //478pi/512
   m_cos[478]  =  14'b11000100000000;     //478pi/512
   m_sin[479]  =  14'b11101010000110;     //479pi/512
   m_cos[479]  =  14'b11000011111000;     //479pi/512
   m_sin[480]  =  14'b11101010011100;     //480pi/512
   m_cos[480]  =  14'b11000011101111;     //480pi/512
   m_sin[481]  =  14'b11101010110011;     //481pi/512
   m_cos[481]  =  14'b11000011100111;     //481pi/512
   m_sin[482]  =  14'b11101011001001;     //482pi/512
   m_cos[482]  =  14'b11000011100000;     //482pi/512
   m_sin[483]  =  14'b11101011100000;     //483pi/512
   m_cos[483]  =  14'b11000011011000;     //483pi/512
   m_sin[484]  =  14'b11101011110110;     //484pi/512
   m_cos[484]  =  14'b11000011010000;     //484pi/512
   m_sin[485]  =  14'b11101100001101;     //485pi/512
   m_cos[485]  =  14'b11000011001001;     //485pi/512
   m_sin[486]  =  14'b11101100100100;     //486pi/512
   m_cos[486]  =  14'b11000011000010;     //486pi/512
   m_sin[487]  =  14'b11101100111011;     //487pi/512
   m_cos[487]  =  14'b11000010111010;     //487pi/512
   m_sin[488]  =  14'b11101101010001;     //488pi/512
   m_cos[488]  =  14'b11000010110011;     //488pi/512
   m_sin[489]  =  14'b11101101101000;     //489pi/512
   m_cos[489]  =  14'b11000010101100;     //489pi/512
   m_sin[490]  =  14'b11101101111111;     //490pi/512
   m_cos[490]  =  14'b11000010100110;     //490pi/512
   m_sin[491]  =  14'b11101110010110;     //491pi/512
   m_cos[491]  =  14'b11000010011111;     //491pi/512
   m_sin[492]  =  14'b11101110101101;     //492pi/512
   m_cos[492]  =  14'b11000010011000;     //492pi/512
   m_sin[493]  =  14'b11101111000100;     //493pi/512
   m_cos[493]  =  14'b11000010010010;     //493pi/512
   m_sin[494]  =  14'b11101111011011;     //494pi/512
   m_cos[494]  =  14'b11000010001100;     //494pi/512
   m_sin[495]  =  14'b11101111110010;     //495pi/512
   m_cos[495]  =  14'b11000010000110;     //495pi/512
   m_sin[496]  =  14'b11110000001001;     //496pi/512
   m_cos[496]  =  14'b11000010000000;     //496pi/512
   m_sin[497]  =  14'b11110000100000;     //497pi/512
   m_cos[497]  =  14'b11000001111010;     //497pi/512
   m_sin[498]  =  14'b11110000111000;     //498pi/512
   m_cos[498]  =  14'b11000001110100;     //498pi/512
   m_sin[499]  =  14'b11110001001111;     //499pi/512
   m_cos[499]  =  14'b11000001101111;     //499pi/512
   m_sin[500]  =  14'b11110001100110;     //500pi/512
   m_cos[500]  =  14'b11000001101001;     //500pi/512
   m_sin[501]  =  14'b11110001111101;     //501pi/512
   m_cos[501]  =  14'b11000001100100;     //501pi/512
   m_sin[502]  =  14'b11110010010101;     //502pi/512
   m_cos[502]  =  14'b11000001011111;     //502pi/512
   m_sin[503]  =  14'b11110010101100;     //503pi/512
   m_cos[503]  =  14'b11000001011010;     //503pi/512
   m_sin[504]  =  14'b11110011000011;     //504pi/512
   m_cos[504]  =  14'b11000001010101;     //504pi/512
   m_sin[505]  =  14'b11110011011011;     //505pi/512
   m_cos[505]  =  14'b11000001010000;     //505pi/512
   m_sin[506]  =  14'b11110011110010;     //506pi/512
   m_cos[506]  =  14'b11000001001011;     //506pi/512
   m_sin[507]  =  14'b11110100001010;     //507pi/512
   m_cos[507]  =  14'b11000001000111;     //507pi/512
   m_sin[508]  =  14'b11110100100001;     //508pi/512
   m_cos[508]  =  14'b11000001000010;     //508pi/512
   m_sin[509]  =  14'b11110100111001;     //509pi/512
   m_cos[509]  =  14'b11000000111110;     //509pi/512
   m_sin[510]  =  14'b11110101010000;     //510pi/512
   m_cos[510]  =  14'b11000000111010;     //510pi/512
   m_sin[511]  =  14'b11110101101000;     //511pi/512
   m_cos[511]  =  14'b11000000110110;     //511pi/512
end

endmodule