module  M_TWIDLE_0_10_v #(parameter stage_FFT = 2, SIZE =10, word_length_tw = 14) (
    input            clk,
    input            en_rd, 
    input   [stage_FFT-2:0]   rd_ptr_angle,

    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );


reg signed [word_length_tw-1:0]  m_cos  [511:0];
reg signed [word_length_tw-1:0]  m_sin  [511:0];

//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd  ) begin
                  cos_data           <= m_cos   [rd_ptr_angle];
                  sin_data           <= m_sin   [rd_ptr_angle];
             end 
        end


//----------------------------------------------------------------------------------------
initial begin


   m_sin[0]  =  14'b00000000000000;     //0pi/512
   m_cos[0]  =  14'b01000000000000;     //0pi/512
   m_sin[1]  =  14'b11111111101001;     //1pi/512
   m_cos[1]  =  14'b00111111111111;     //1pi/512
   m_sin[2]  =  14'b11111111010011;     //2pi/512
   m_cos[2]  =  14'b00111111111111;     //2pi/512
   m_sin[3]  =  14'b11111110111100;     //3pi/512
   m_cos[3]  =  14'b00111111111111;     //3pi/512
   m_sin[4]  =  14'b11111110100110;     //4pi/512
   m_cos[4]  =  14'b00111111111111;     //4pi/512
   m_sin[5]  =  14'b11111110001111;     //5pi/512
   m_cos[5]  =  14'b00111111111110;     //5pi/512
   m_sin[6]  =  14'b11111101111000;     //6pi/512
   m_cos[6]  =  14'b00111111111101;     //6pi/512
   m_sin[7]  =  14'b11111101100010;     //7pi/512
   m_cos[7]  =  14'b00111111111100;     //7pi/512
   m_sin[8]  =  14'b11111101001011;     //8pi/512
   m_cos[8]  =  14'b00111111111100;     //8pi/512
   m_sin[9]  =  14'b11111100110101;     //9pi/512
   m_cos[9]  =  14'b00111111111010;     //9pi/512
   m_sin[10]  =  14'b11111100011110;     //10pi/512
   m_cos[10]  =  14'b00111111111001;     //10pi/512
   m_sin[11]  =  14'b11111100000111;     //11pi/512
   m_cos[11]  =  14'b00111111111000;     //11pi/512
   m_sin[12]  =  14'b11111011110001;     //12pi/512
   m_cos[12]  =  14'b00111111110111;     //12pi/512
   m_sin[13]  =  14'b11111011011010;     //13pi/512
   m_cos[13]  =  14'b00111111110101;     //13pi/512
   m_sin[14]  =  14'b11111011000100;     //14pi/512
   m_cos[14]  =  14'b00111111110011;     //14pi/512
   m_sin[15]  =  14'b11111010101101;     //15pi/512
   m_cos[15]  =  14'b00111111110001;     //15pi/512
   m_sin[16]  =  14'b11111010010111;     //16pi/512
   m_cos[16]  =  14'b00111111110000;     //16pi/512
   m_sin[17]  =  14'b11111010000000;     //17pi/512
   m_cos[17]  =  14'b00111111101101;     //17pi/512
   m_sin[18]  =  14'b11111001101010;     //18pi/512
   m_cos[18]  =  14'b00111111101011;     //18pi/512
   m_sin[19]  =  14'b11111001010011;     //19pi/512
   m_cos[19]  =  14'b00111111101001;     //19pi/512
   m_sin[20]  =  14'b11111000111101;     //20pi/512
   m_cos[20]  =  14'b00111111100111;     //20pi/512
   m_sin[21]  =  14'b11111000100110;     //21pi/512
   m_cos[21]  =  14'b00111111100100;     //21pi/512
   m_sin[22]  =  14'b11111000010000;     //22pi/512
   m_cos[22]  =  14'b00111111100001;     //22pi/512
   m_sin[23]  =  14'b11110111111001;     //23pi/512
   m_cos[23]  =  14'b00111111011111;     //23pi/512
   m_sin[24]  =  14'b11110111100011;     //24pi/512
   m_cos[24]  =  14'b00111111011100;     //24pi/512
   m_sin[25]  =  14'b11110111001100;     //25pi/512
   m_cos[25]  =  14'b00111111011001;     //25pi/512
   m_sin[26]  =  14'b11110110110110;     //26pi/512
   m_cos[26]  =  14'b00111111010101;     //26pi/512
   m_sin[27]  =  14'b11110110100000;     //27pi/512
   m_cos[27]  =  14'b00111111010010;     //27pi/512
   m_sin[28]  =  14'b11110110001001;     //28pi/512
   m_cos[28]  =  14'b00111111001111;     //28pi/512
   m_sin[29]  =  14'b11110101110011;     //29pi/512
   m_cos[29]  =  14'b00111111001011;     //29pi/512
   m_sin[30]  =  14'b11110101011101;     //30pi/512
   m_cos[30]  =  14'b00111111000111;     //30pi/512
   m_sin[31]  =  14'b11110101000110;     //31pi/512
   m_cos[31]  =  14'b00111111000100;     //31pi/512
   m_sin[32]  =  14'b11110100110000;     //32pi/512
   m_cos[32]  =  14'b00111111000000;     //32pi/512
   m_sin[33]  =  14'b11110100011010;     //33pi/512
   m_cos[33]  =  14'b00111110111100;     //33pi/512
   m_sin[34]  =  14'b11110100000011;     //34pi/512
   m_cos[34]  =  14'b00111110111000;     //34pi/512
   m_sin[35]  =  14'b11110011101101;     //35pi/512
   m_cos[35]  =  14'b00111110110011;     //35pi/512
   m_sin[36]  =  14'b11110011010111;     //36pi/512
   m_cos[36]  =  14'b00111110101111;     //36pi/512
   m_sin[37]  =  14'b11110011000001;     //37pi/512
   m_cos[37]  =  14'b00111110101010;     //37pi/512
   m_sin[38]  =  14'b11110010101011;     //38pi/512
   m_cos[38]  =  14'b00111110100110;     //38pi/512
   m_sin[39]  =  14'b11110010010101;     //39pi/512
   m_cos[39]  =  14'b00111110100001;     //39pi/512
   m_sin[40]  =  14'b11110001111111;     //40pi/512
   m_cos[40]  =  14'b00111110011100;     //40pi/512
   m_sin[41]  =  14'b11110001101001;     //41pi/512
   m_cos[41]  =  14'b00111110010111;     //41pi/512
   m_sin[42]  =  14'b11110001010010;     //42pi/512
   m_cos[42]  =  14'b00111110010010;     //42pi/512
   m_sin[43]  =  14'b11110000111100;     //43pi/512
   m_cos[43]  =  14'b00111110001101;     //43pi/512
   m_sin[44]  =  14'b11110000100111;     //44pi/512
   m_cos[44]  =  14'b00111110000111;     //44pi/512
   m_sin[45]  =  14'b11110000010001;     //45pi/512
   m_cos[45]  =  14'b00111110000010;     //45pi/512
   m_sin[46]  =  14'b11101111111011;     //46pi/512
   m_cos[46]  =  14'b00111101111100;     //46pi/512
   m_sin[47]  =  14'b11101111100101;     //47pi/512
   m_cos[47]  =  14'b00111101110110;     //47pi/512
   m_sin[48]  =  14'b11101111001111;     //48pi/512
   m_cos[48]  =  14'b00111101110000;     //48pi/512
   m_sin[49]  =  14'b11101110111001;     //49pi/512
   m_cos[49]  =  14'b00111101101010;     //49pi/512
   m_sin[50]  =  14'b11101110100011;     //50pi/512
   m_cos[50]  =  14'b00111101100100;     //50pi/512
   m_sin[51]  =  14'b11101110001110;     //51pi/512
   m_cos[51]  =  14'b00111101011110;     //51pi/512
   m_sin[52]  =  14'b11101101111000;     //52pi/512
   m_cos[52]  =  14'b00111101011000;     //52pi/512
   m_sin[53]  =  14'b11101101100010;     //53pi/512
   m_cos[53]  =  14'b00111101010001;     //53pi/512
   m_sin[54]  =  14'b11101101001101;     //54pi/512
   m_cos[54]  =  14'b00111101001011;     //54pi/512
   m_sin[55]  =  14'b11101100110111;     //55pi/512
   m_cos[55]  =  14'b00111101000100;     //55pi/512
   m_sin[56]  =  14'b11101100100001;     //56pi/512
   m_cos[56]  =  14'b00111100111101;     //56pi/512
   m_sin[57]  =  14'b11101100001100;     //57pi/512
   m_cos[57]  =  14'b00111100110110;     //57pi/512
   m_sin[58]  =  14'b11101011110110;     //58pi/512
   m_cos[58]  =  14'b00111100101111;     //58pi/512
   m_sin[59]  =  14'b11101011100001;     //59pi/512
   m_cos[59]  =  14'b00111100101000;     //59pi/512
   m_sin[60]  =  14'b11101011001100;     //60pi/512
   m_cos[60]  =  14'b00111100100001;     //60pi/512
   m_sin[61]  =  14'b11101010110110;     //61pi/512
   m_cos[61]  =  14'b00111100011001;     //61pi/512
   m_sin[62]  =  14'b11101010100001;     //62pi/512
   m_cos[62]  =  14'b00111100010010;     //62pi/512
   m_sin[63]  =  14'b11101010001100;     //63pi/512
   m_cos[63]  =  14'b00111100001010;     //63pi/512
   m_sin[64]  =  14'b11101001110110;     //64pi/512
   m_cos[64]  =  14'b00111100000010;     //64pi/512
   m_sin[65]  =  14'b11101001100001;     //65pi/512
   m_cos[65]  =  14'b00111011111010;     //65pi/512
   m_sin[66]  =  14'b11101001001100;     //66pi/512
   m_cos[66]  =  14'b00111011110010;     //66pi/512
   m_sin[67]  =  14'b11101000110111;     //67pi/512
   m_cos[67]  =  14'b00111011101010;     //67pi/512
   m_sin[68]  =  14'b11101000100010;     //68pi/512
   m_cos[68]  =  14'b00111011100010;     //68pi/512
   m_sin[69]  =  14'b11101000001101;     //69pi/512
   m_cos[69]  =  14'b00111011011010;     //69pi/512
   m_sin[70]  =  14'b11100111111000;     //70pi/512
   m_cos[70]  =  14'b00111011010001;     //70pi/512
   m_sin[71]  =  14'b11100111100011;     //71pi/512
   m_cos[71]  =  14'b00111011001001;     //71pi/512
   m_sin[72]  =  14'b11100111001110;     //72pi/512
   m_cos[72]  =  14'b00111011000000;     //72pi/512
   m_sin[73]  =  14'b11100110111001;     //73pi/512
   m_cos[73]  =  14'b00111010110111;     //73pi/512
   m_sin[74]  =  14'b11100110100100;     //74pi/512
   m_cos[74]  =  14'b00111010101110;     //74pi/512
   m_sin[75]  =  14'b11100110010000;     //75pi/512
   m_cos[75]  =  14'b00111010100101;     //75pi/512
   m_sin[76]  =  14'b11100101111011;     //76pi/512
   m_cos[76]  =  14'b00111010011100;     //76pi/512
   m_sin[77]  =  14'b11100101100110;     //77pi/512
   m_cos[77]  =  14'b00111010010011;     //77pi/512
   m_sin[78]  =  14'b11100101010010;     //78pi/512
   m_cos[78]  =  14'b00111010001001;     //78pi/512
   m_sin[79]  =  14'b11100100111101;     //79pi/512
   m_cos[79]  =  14'b00111010000000;     //79pi/512
   m_sin[80]  =  14'b11100100101001;     //80pi/512
   m_cos[80]  =  14'b00111001110110;     //80pi/512
   m_sin[81]  =  14'b11100100010100;     //81pi/512
   m_cos[81]  =  14'b00111001101101;     //81pi/512
   m_sin[82]  =  14'b11100100000000;     //82pi/512
   m_cos[82]  =  14'b00111001100011;     //82pi/512
   m_sin[83]  =  14'b11100011101100;     //83pi/512
   m_cos[83]  =  14'b00111001011001;     //83pi/512
   m_sin[84]  =  14'b11100011010111;     //84pi/512
   m_cos[84]  =  14'b00111001001111;     //84pi/512
   m_sin[85]  =  14'b11100011000011;     //85pi/512
   m_cos[85]  =  14'b00111001000100;     //85pi/512
   m_sin[86]  =  14'b11100010101111;     //86pi/512
   m_cos[86]  =  14'b00111000111010;     //86pi/512
   m_sin[87]  =  14'b11100010011011;     //87pi/512
   m_cos[87]  =  14'b00111000110000;     //87pi/512
   m_sin[88]  =  14'b11100010000111;     //88pi/512
   m_cos[88]  =  14'b00111000100101;     //88pi/512
   m_sin[89]  =  14'b11100001110011;     //89pi/512
   m_cos[89]  =  14'b00111000011011;     //89pi/512
   m_sin[90]  =  14'b11100001011111;     //90pi/512
   m_cos[90]  =  14'b00111000010000;     //90pi/512
   m_sin[91]  =  14'b11100001001011;     //91pi/512
   m_cos[91]  =  14'b00111000000101;     //91pi/512
   m_sin[92]  =  14'b11100000110111;     //92pi/512
   m_cos[92]  =  14'b00110111111010;     //92pi/512
   m_sin[93]  =  14'b11100000100100;     //93pi/512
   m_cos[93]  =  14'b00110111101111;     //93pi/512
   m_sin[94]  =  14'b11100000010000;     //94pi/512
   m_cos[94]  =  14'b00110111100100;     //94pi/512
   m_sin[95]  =  14'b11011111111100;     //95pi/512
   m_cos[95]  =  14'b00110111011001;     //95pi/512
   m_sin[96]  =  14'b11011111101001;     //96pi/512
   m_cos[96]  =  14'b00110111001101;     //96pi/512
   m_sin[97]  =  14'b11011111010101;     //97pi/512
   m_cos[97]  =  14'b00110111000010;     //97pi/512
   m_sin[98]  =  14'b11011111000010;     //98pi/512
   m_cos[98]  =  14'b00110110110110;     //98pi/512
   m_sin[99]  =  14'b11011110101111;     //99pi/512
   m_cos[99]  =  14'b00110110101010;     //99pi/512
   m_sin[100]  =  14'b11011110011011;     //100pi/512
   m_cos[100]  =  14'b00110110011111;     //100pi/512
   m_sin[101]  =  14'b11011110001000;     //101pi/512
   m_cos[101]  =  14'b00110110010011;     //101pi/512
   m_sin[102]  =  14'b11011101110101;     //102pi/512
   m_cos[102]  =  14'b00110110000111;     //102pi/512
   m_sin[103]  =  14'b11011101100010;     //103pi/512
   m_cos[103]  =  14'b00110101111011;     //103pi/512
   m_sin[104]  =  14'b11011101001111;     //104pi/512
   m_cos[104]  =  14'b00110101101110;     //104pi/512
   m_sin[105]  =  14'b11011100111100;     //105pi/512
   m_cos[105]  =  14'b00110101100010;     //105pi/512
   m_sin[106]  =  14'b11011100101001;     //106pi/512
   m_cos[106]  =  14'b00110101010110;     //106pi/512
   m_sin[107]  =  14'b11011100010110;     //107pi/512
   m_cos[107]  =  14'b00110101001001;     //107pi/512
   m_sin[108]  =  14'b11011100000011;     //108pi/512
   m_cos[108]  =  14'b00110100111100;     //108pi/512
   m_sin[109]  =  14'b11011011110001;     //109pi/512
   m_cos[109]  =  14'b00110100110000;     //109pi/512
   m_sin[110]  =  14'b11011011011110;     //110pi/512
   m_cos[110]  =  14'b00110100100011;     //110pi/512
   m_sin[111]  =  14'b11011011001100;     //111pi/512
   m_cos[111]  =  14'b00110100010110;     //111pi/512
   m_sin[112]  =  14'b11011010111001;     //112pi/512
   m_cos[112]  =  14'b00110100001001;     //112pi/512
   m_sin[113]  =  14'b11011010100111;     //113pi/512
   m_cos[113]  =  14'b00110011111100;     //113pi/512
   m_sin[114]  =  14'b11011010010100;     //114pi/512
   m_cos[114]  =  14'b00110011101110;     //114pi/512
   m_sin[115]  =  14'b11011010000010;     //115pi/512
   m_cos[115]  =  14'b00110011100001;     //115pi/512
   m_sin[116]  =  14'b11011001110000;     //116pi/512
   m_cos[116]  =  14'b00110011010011;     //116pi/512
   m_sin[117]  =  14'b11011001011110;     //117pi/512
   m_cos[117]  =  14'b00110011000110;     //117pi/512
   m_sin[118]  =  14'b11011001001100;     //118pi/512
   m_cos[118]  =  14'b00110010111000;     //118pi/512
   m_sin[119]  =  14'b11011000111010;     //119pi/512
   m_cos[119]  =  14'b00110010101010;     //119pi/512
   m_sin[120]  =  14'b11011000101000;     //120pi/512
   m_cos[120]  =  14'b00110010011101;     //120pi/512
   m_sin[121]  =  14'b11011000010110;     //121pi/512
   m_cos[121]  =  14'b00110010001111;     //121pi/512
   m_sin[122]  =  14'b11011000000101;     //122pi/512
   m_cos[122]  =  14'b00110010000001;     //122pi/512
   m_sin[123]  =  14'b11010111110011;     //123pi/512
   m_cos[123]  =  14'b00110001110010;     //123pi/512
   m_sin[124]  =  14'b11010111100001;     //124pi/512
   m_cos[124]  =  14'b00110001100100;     //124pi/512
   m_sin[125]  =  14'b11010111010000;     //125pi/512
   m_cos[125]  =  14'b00110001010110;     //125pi/512
   m_sin[126]  =  14'b11010110111110;     //126pi/512
   m_cos[126]  =  14'b00110001000111;     //126pi/512
   m_sin[127]  =  14'b11010110101101;     //127pi/512
   m_cos[127]  =  14'b00110000111001;     //127pi/512
   m_sin[128]  =  14'b11010110011100;     //128pi/512
   m_cos[128]  =  14'b00110000101010;     //128pi/512
   m_sin[129]  =  14'b11010110001011;     //129pi/512
   m_cos[129]  =  14'b00110000011011;     //129pi/512
   m_sin[130]  =  14'b11010101111010;     //130pi/512
   m_cos[130]  =  14'b00110000001101;     //130pi/512
   m_sin[131]  =  14'b11010101101001;     //131pi/512
   m_cos[131]  =  14'b00101111111110;     //131pi/512
   m_sin[132]  =  14'b11010101011000;     //132pi/512
   m_cos[132]  =  14'b00101111101111;     //132pi/512
   m_sin[133]  =  14'b11010101000111;     //133pi/512
   m_cos[133]  =  14'b00101111011111;     //133pi/512
   m_sin[134]  =  14'b11010100110110;     //134pi/512
   m_cos[134]  =  14'b00101111010000;     //134pi/512
   m_sin[135]  =  14'b11010100100101;     //135pi/512
   m_cos[135]  =  14'b00101111000001;     //135pi/512
   m_sin[136]  =  14'b11010100010101;     //136pi/512
   m_cos[136]  =  14'b00101110110010;     //136pi/512
   m_sin[137]  =  14'b11010100000100;     //137pi/512
   m_cos[137]  =  14'b00101110100010;     //137pi/512
   m_sin[138]  =  14'b11010011110100;     //138pi/512
   m_cos[138]  =  14'b00101110010011;     //138pi/512
   m_sin[139]  =  14'b11010011100100;     //139pi/512
   m_cos[139]  =  14'b00101110000011;     //139pi/512
   m_sin[140]  =  14'b11010011010011;     //140pi/512
   m_cos[140]  =  14'b00101101110011;     //140pi/512
   m_sin[141]  =  14'b11010011000011;     //141pi/512
   m_cos[141]  =  14'b00101101100011;     //141pi/512
   m_sin[142]  =  14'b11010010110011;     //142pi/512
   m_cos[142]  =  14'b00101101010011;     //142pi/512
   m_sin[143]  =  14'b11010010100011;     //143pi/512
   m_cos[143]  =  14'b00101101000011;     //143pi/512
   m_sin[144]  =  14'b11010010010011;     //144pi/512
   m_cos[144]  =  14'b00101100110011;     //144pi/512
   m_sin[145]  =  14'b11010010000100;     //145pi/512
   m_cos[145]  =  14'b00101100100011;     //145pi/512
   m_sin[146]  =  14'b11010001110100;     //146pi/512
   m_cos[146]  =  14'b00101100010011;     //146pi/512
   m_sin[147]  =  14'b11010001100100;     //147pi/512
   m_cos[147]  =  14'b00101100000010;     //147pi/512
   m_sin[148]  =  14'b11010001010101;     //148pi/512
   m_cos[148]  =  14'b00101011110010;     //148pi/512
   m_sin[149]  =  14'b11010001000101;     //149pi/512
   m_cos[149]  =  14'b00101011100001;     //149pi/512
   m_sin[150]  =  14'b11010000110110;     //150pi/512
   m_cos[150]  =  14'b00101011010001;     //150pi/512
   m_sin[151]  =  14'b11010000100111;     //151pi/512
   m_cos[151]  =  14'b00101011000000;     //151pi/512
   m_sin[152]  =  14'b11010000011000;     //152pi/512
   m_cos[152]  =  14'b00101010101111;     //152pi/512
   m_sin[153]  =  14'b11010000001001;     //153pi/512
   m_cos[153]  =  14'b00101010011110;     //153pi/512
   m_sin[154]  =  14'b11001111111010;     //154pi/512
   m_cos[154]  =  14'b00101010001101;     //154pi/512
   m_sin[155]  =  14'b11001111101011;     //155pi/512
   m_cos[155]  =  14'b00101001111100;     //155pi/512
   m_sin[156]  =  14'b11001111011100;     //156pi/512
   m_cos[156]  =  14'b00101001101011;     //156pi/512
   m_sin[157]  =  14'b11001111001101;     //157pi/512
   m_cos[157]  =  14'b00101001011010;     //157pi/512
   m_sin[158]  =  14'b11001110111111;     //158pi/512
   m_cos[158]  =  14'b00101001001001;     //158pi/512
   m_sin[159]  =  14'b11001110110000;     //159pi/512
   m_cos[159]  =  14'b00101000110111;     //159pi/512
   m_sin[160]  =  14'b11001110100010;     //160pi/512
   m_cos[160]  =  14'b00101000100110;     //160pi/512
   m_sin[161]  =  14'b11001110010011;     //161pi/512
   m_cos[161]  =  14'b00101000010100;     //161pi/512
   m_sin[162]  =  14'b11001110000101;     //162pi/512
   m_cos[162]  =  14'b00101000000011;     //162pi/512
   m_sin[163]  =  14'b11001101110111;     //163pi/512
   m_cos[163]  =  14'b00100111110001;     //163pi/512
   m_sin[164]  =  14'b11001101101001;     //164pi/512
   m_cos[164]  =  14'b00100111011111;     //164pi/512
   m_sin[165]  =  14'b11001101011011;     //165pi/512
   m_cos[165]  =  14'b00100111001110;     //165pi/512
   m_sin[166]  =  14'b11001101001101;     //166pi/512
   m_cos[166]  =  14'b00100110111100;     //166pi/512
   m_sin[167]  =  14'b11001101000000;     //167pi/512
   m_cos[167]  =  14'b00100110101010;     //167pi/512
   m_sin[168]  =  14'b11001100110010;     //168pi/512
   m_cos[168]  =  14'b00100110011000;     //168pi/512
   m_sin[169]  =  14'b11001100100101;     //169pi/512
   m_cos[169]  =  14'b00100110000101;     //169pi/512
   m_sin[170]  =  14'b11001100010111;     //170pi/512
   m_cos[170]  =  14'b00100101110011;     //170pi/512
   m_sin[171]  =  14'b11001100001010;     //171pi/512
   m_cos[171]  =  14'b00100101100001;     //171pi/512
   m_sin[172]  =  14'b11001011111101;     //172pi/512
   m_cos[172]  =  14'b00100101001111;     //172pi/512
   m_sin[173]  =  14'b11001011110000;     //173pi/512
   m_cos[173]  =  14'b00100100111100;     //173pi/512
   m_sin[174]  =  14'b11001011100011;     //174pi/512
   m_cos[174]  =  14'b00100100101010;     //174pi/512
   m_sin[175]  =  14'b11001011010110;     //175pi/512
   m_cos[175]  =  14'b00100100010111;     //175pi/512
   m_sin[176]  =  14'b11001011001001;     //176pi/512
   m_cos[176]  =  14'b00100100000100;     //176pi/512
   m_sin[177]  =  14'b11001010111100;     //177pi/512
   m_cos[177]  =  14'b00100011110010;     //177pi/512
   m_sin[178]  =  14'b11001010110000;     //178pi/512
   m_cos[178]  =  14'b00100011011111;     //178pi/512
   m_sin[179]  =  14'b11001010100011;     //179pi/512
   m_cos[179]  =  14'b00100011001100;     //179pi/512
   m_sin[180]  =  14'b11001010010111;     //180pi/512
   m_cos[180]  =  14'b00100010111001;     //180pi/512
   m_sin[181]  =  14'b11001010001010;     //181pi/512
   m_cos[181]  =  14'b00100010100110;     //181pi/512
   m_sin[182]  =  14'b11001001111110;     //182pi/512
   m_cos[182]  =  14'b00100010010011;     //182pi/512
   m_sin[183]  =  14'b11001001110010;     //183pi/512
   m_cos[183]  =  14'b00100010000000;     //183pi/512
   m_sin[184]  =  14'b11001001100110;     //184pi/512
   m_cos[184]  =  14'b00100001101101;     //184pi/512
   m_sin[185]  =  14'b11001001011010;     //185pi/512
   m_cos[185]  =  14'b00100001011010;     //185pi/512
   m_sin[186]  =  14'b11001001001111;     //186pi/512
   m_cos[186]  =  14'b00100001000110;     //186pi/512
   m_sin[187]  =  14'b11001001000011;     //187pi/512
   m_cos[187]  =  14'b00100000110011;     //187pi/512
   m_sin[188]  =  14'b11001000110111;     //188pi/512
   m_cos[188]  =  14'b00100000011111;     //188pi/512
   m_sin[189]  =  14'b11001000101100;     //189pi/512
   m_cos[189]  =  14'b00100000001100;     //189pi/512
   m_sin[190]  =  14'b11001000100001;     //190pi/512
   m_cos[190]  =  14'b00011111111000;     //190pi/512
   m_sin[191]  =  14'b11001000010101;     //191pi/512
   m_cos[191]  =  14'b00011111100101;     //191pi/512
   m_sin[192]  =  14'b11001000001010;     //192pi/512
   m_cos[192]  =  14'b00011111010001;     //192pi/512
   m_sin[193]  =  14'b11000111111111;     //193pi/512
   m_cos[193]  =  14'b00011110111101;     //193pi/512
   m_sin[194]  =  14'b11000111110100;     //194pi/512
   m_cos[194]  =  14'b00011110101001;     //194pi/512
   m_sin[195]  =  14'b11000111101010;     //195pi/512
   m_cos[195]  =  14'b00011110010101;     //195pi/512
   m_sin[196]  =  14'b11000111011111;     //196pi/512
   m_cos[196]  =  14'b00011110000001;     //196pi/512
   m_sin[197]  =  14'b11000111010100;     //197pi/512
   m_cos[197]  =  14'b00011101101101;     //197pi/512
   m_sin[198]  =  14'b11000111001010;     //198pi/512
   m_cos[198]  =  14'b00011101011001;     //198pi/512
   m_sin[199]  =  14'b11000111000000;     //199pi/512
   m_cos[199]  =  14'b00011101000101;     //199pi/512
   m_sin[200]  =  14'b11000110110101;     //200pi/512
   m_cos[200]  =  14'b00011100110001;     //200pi/512
   m_sin[201]  =  14'b11000110101011;     //201pi/512
   m_cos[201]  =  14'b00011100011101;     //201pi/512
   m_sin[202]  =  14'b11000110100001;     //202pi/512
   m_cos[202]  =  14'b00011100001001;     //202pi/512
   m_sin[203]  =  14'b11000110010111;     //203pi/512
   m_cos[203]  =  14'b00011011110100;     //203pi/512
   m_sin[204]  =  14'b11000110001110;     //204pi/512
   m_cos[204]  =  14'b00011011100000;     //204pi/512
   m_sin[205]  =  14'b11000110000100;     //205pi/512
   m_cos[205]  =  14'b00011011001011;     //205pi/512
   m_sin[206]  =  14'b11000101111010;     //206pi/512
   m_cos[206]  =  14'b00011010110111;     //206pi/512
   m_sin[207]  =  14'b11000101110001;     //207pi/512
   m_cos[207]  =  14'b00011010100010;     //207pi/512
   m_sin[208]  =  14'b11000101101000;     //208pi/512
   m_cos[208]  =  14'b00011010001110;     //208pi/512
   m_sin[209]  =  14'b11000101011110;     //209pi/512
   m_cos[209]  =  14'b00011001111001;     //209pi/512
   m_sin[210]  =  14'b11000101010101;     //210pi/512
   m_cos[210]  =  14'b00011001100100;     //210pi/512
   m_sin[211]  =  14'b11000101001100;     //211pi/512
   m_cos[211]  =  14'b00011001010000;     //211pi/512
   m_sin[212]  =  14'b11000101000011;     //212pi/512
   m_cos[212]  =  14'b00011000111011;     //212pi/512
   m_sin[213]  =  14'b11000100111011;     //213pi/512
   m_cos[213]  =  14'b00011000100110;     //213pi/512
   m_sin[214]  =  14'b11000100110010;     //214pi/512
   m_cos[214]  =  14'b00011000010001;     //214pi/512
   m_sin[215]  =  14'b11000100101010;     //215pi/512
   m_cos[215]  =  14'b00010111111100;     //215pi/512
   m_sin[216]  =  14'b11000100100001;     //216pi/512
   m_cos[216]  =  14'b00010111100111;     //216pi/512
   m_sin[217]  =  14'b11000100011001;     //217pi/512
   m_cos[217]  =  14'b00010111010010;     //217pi/512
   m_sin[218]  =  14'b11000100010001;     //218pi/512
   m_cos[218]  =  14'b00010110111101;     //218pi/512
   m_sin[219]  =  14'b11000100001001;     //219pi/512
   m_cos[219]  =  14'b00010110101000;     //219pi/512
   m_sin[220]  =  14'b11000100000001;     //220pi/512
   m_cos[220]  =  14'b00010110010011;     //220pi/512
   m_sin[221]  =  14'b11000011111001;     //221pi/512
   m_cos[221]  =  14'b00010101111101;     //221pi/512
   m_sin[222]  =  14'b11000011110001;     //222pi/512
   m_cos[222]  =  14'b00010101101000;     //222pi/512
   m_sin[223]  =  14'b11000011101010;     //223pi/512
   m_cos[223]  =  14'b00010101010011;     //223pi/512
   m_sin[224]  =  14'b11000011100010;     //224pi/512
   m_cos[224]  =  14'b00010100111101;     //224pi/512
   m_sin[225]  =  14'b11000011011011;     //225pi/512
   m_cos[225]  =  14'b00010100101000;     //225pi/512
   m_sin[226]  =  14'b11000011010011;     //226pi/512
   m_cos[226]  =  14'b00010100010011;     //226pi/512
   m_sin[227]  =  14'b11000011001100;     //227pi/512
   m_cos[227]  =  14'b00010011111101;     //227pi/512
   m_sin[228]  =  14'b11000011000101;     //228pi/512
   m_cos[228]  =  14'b00010011101000;     //228pi/512
   m_sin[229]  =  14'b11000010111111;     //229pi/512
   m_cos[229]  =  14'b00010011010010;     //229pi/512
   m_sin[230]  =  14'b11000010111000;     //230pi/512
   m_cos[230]  =  14'b00010010111101;     //230pi/512
   m_sin[231]  =  14'b11000010110001;     //231pi/512
   m_cos[231]  =  14'b00010010100111;     //231pi/512
   m_sin[232]  =  14'b11000010101011;     //232pi/512
   m_cos[232]  =  14'b00010010010001;     //232pi/512
   m_sin[233]  =  14'b11000010100100;     //233pi/512
   m_cos[233]  =  14'b00010001111100;     //233pi/512
   m_sin[234]  =  14'b11000010011110;     //234pi/512
   m_cos[234]  =  14'b00010001100110;     //234pi/512
   m_sin[235]  =  14'b11000010011000;     //235pi/512
   m_cos[235]  =  14'b00010001010000;     //235pi/512
   m_sin[236]  =  14'b11000010010010;     //236pi/512
   m_cos[236]  =  14'b00010000111010;     //236pi/512
   m_sin[237]  =  14'b11000010001100;     //237pi/512
   m_cos[237]  =  14'b00010000100100;     //237pi/512
   m_sin[238]  =  14'b11000010000110;     //238pi/512
   m_cos[238]  =  14'b00010000001111;     //238pi/512
   m_sin[239]  =  14'b11000010000000;     //239pi/512
   m_cos[239]  =  14'b00001111111001;     //239pi/512
   m_sin[240]  =  14'b11000001111011;     //240pi/512
   m_cos[240]  =  14'b00001111100011;     //240pi/512
   m_sin[241]  =  14'b11000001110101;     //241pi/512
   m_cos[241]  =  14'b00001111001101;     //241pi/512
   m_sin[242]  =  14'b11000001110000;     //242pi/512
   m_cos[242]  =  14'b00001110110111;     //242pi/512
   m_sin[243]  =  14'b11000001101011;     //243pi/512
   m_cos[243]  =  14'b00001110100001;     //243pi/512
   m_sin[244]  =  14'b11000001100110;     //244pi/512
   m_cos[244]  =  14'b00001110001011;     //244pi/512
   m_sin[245]  =  14'b11000001100001;     //245pi/512
   m_cos[245]  =  14'b00001101110101;     //245pi/512
   m_sin[246]  =  14'b11000001011100;     //246pi/512
   m_cos[246]  =  14'b00001101011111;     //246pi/512
   m_sin[247]  =  14'b11000001010111;     //247pi/512
   m_cos[247]  =  14'b00001101001000;     //247pi/512
   m_sin[248]  =  14'b11000001010011;     //248pi/512
   m_cos[248]  =  14'b00001100110010;     //248pi/512
   m_sin[249]  =  14'b11000001001110;     //249pi/512
   m_cos[249]  =  14'b00001100011100;     //249pi/512
   m_sin[250]  =  14'b11000001001010;     //250pi/512
   m_cos[250]  =  14'b00001100000110;     //250pi/512
   m_sin[251]  =  14'b11000001000110;     //251pi/512
   m_cos[251]  =  14'b00001011110000;     //251pi/512
   m_sin[252]  =  14'b11000001000010;     //252pi/512
   m_cos[252]  =  14'b00001011011001;     //252pi/512
   m_sin[253]  =  14'b11000000111110;     //253pi/512
   m_cos[253]  =  14'b00001011000011;     //253pi/512
   m_sin[254]  =  14'b11000000111010;     //254pi/512
   m_cos[254]  =  14'b00001010101101;     //254pi/512
   m_sin[255]  =  14'b11000000110110;     //255pi/512
   m_cos[255]  =  14'b00001010010111;     //255pi/512
   m_sin[256]  =  14'b11000000110010;     //256pi/512
   m_cos[256]  =  14'b00001010000000;     //256pi/512
   m_sin[257]  =  14'b11000000101111;     //257pi/512
   m_cos[257]  =  14'b00001001101010;     //257pi/512
   m_sin[258]  =  14'b11000000101100;     //258pi/512
   m_cos[258]  =  14'b00001001010100;     //258pi/512
   m_sin[259]  =  14'b11000000101000;     //259pi/512
   m_cos[259]  =  14'b00001000111101;     //259pi/512
   m_sin[260]  =  14'b11000000100101;     //260pi/512
   m_cos[260]  =  14'b00001000100111;     //260pi/512
   m_sin[261]  =  14'b11000000100010;     //261pi/512
   m_cos[261]  =  14'b00001000010000;     //261pi/512
   m_sin[262]  =  14'b11000000011111;     //262pi/512
   m_cos[262]  =  14'b00000111111010;     //262pi/512
   m_sin[263]  =  14'b11000000011101;     //263pi/512
   m_cos[263]  =  14'b00000111100011;     //263pi/512
   m_sin[264]  =  14'b11000000011010;     //264pi/512
   m_cos[264]  =  14'b00000111001101;     //264pi/512
   m_sin[265]  =  14'b11000000011000;     //265pi/512
   m_cos[265]  =  14'b00000110110110;     //265pi/512
   m_sin[266]  =  14'b11000000010101;     //266pi/512
   m_cos[266]  =  14'b00000110100000;     //266pi/512
   m_sin[267]  =  14'b11000000010011;     //267pi/512
   m_cos[267]  =  14'b00000110001001;     //267pi/512
   m_sin[268]  =  14'b11000000010001;     //268pi/512
   m_cos[268]  =  14'b00000101110011;     //268pi/512
   m_sin[269]  =  14'b11000000001111;     //269pi/512
   m_cos[269]  =  14'b00000101011100;     //269pi/512
   m_sin[270]  =  14'b11000000001101;     //270pi/512
   m_cos[270]  =  14'b00000101000110;     //270pi/512
   m_sin[271]  =  14'b11000000001011;     //271pi/512
   m_cos[271]  =  14'b00000100101111;     //271pi/512
   m_sin[272]  =  14'b11000000001010;     //272pi/512
   m_cos[272]  =  14'b00000100011001;     //272pi/512
   m_sin[273]  =  14'b11000000001000;     //273pi/512
   m_cos[273]  =  14'b00000100000010;     //273pi/512
   m_sin[274]  =  14'b11000000000111;     //274pi/512
   m_cos[274]  =  14'b00000011101100;     //274pi/512
   m_sin[275]  =  14'b11000000000110;     //275pi/512
   m_cos[275]  =  14'b00000011010101;     //275pi/512
   m_sin[276]  =  14'b11000000000100;     //276pi/512
   m_cos[276]  =  14'b00000010111110;     //276pi/512
   m_sin[277]  =  14'b11000000000011;     //277pi/512
   m_cos[277]  =  14'b00000010101000;     //277pi/512
   m_sin[278]  =  14'b11000000000011;     //278pi/512
   m_cos[278]  =  14'b00000010010001;     //278pi/512
   m_sin[279]  =  14'b11000000000010;     //279pi/512
   m_cos[279]  =  14'b00000001111011;     //279pi/512
   m_sin[280]  =  14'b11000000000001;     //280pi/512
   m_cos[280]  =  14'b00000001100100;     //280pi/512
   m_sin[281]  =  14'b11000000000001;     //281pi/512
   m_cos[281]  =  14'b00000001001101;     //281pi/512
   m_sin[282]  =  14'b11000000000000;     //282pi/512
   m_cos[282]  =  14'b00000000110111;     //282pi/512
   m_sin[283]  =  14'b11000000000000;     //283pi/512
   m_cos[283]  =  14'b00000000100000;     //283pi/512
   m_sin[284]  =  14'b11000000000000;     //284pi/512
   m_cos[284]  =  14'b00000000001010;     //284pi/512
   m_sin[285]  =  14'b11000000000000;     //285pi/512
   m_cos[285]  =  14'b11111111110011;     //285pi/512
   m_sin[286]  =  14'b11000000000000;     //286pi/512
   m_cos[286]  =  14'b11111111011101;     //286pi/512
   m_sin[287]  =  14'b11000000000000;     //287pi/512
   m_cos[287]  =  14'b11111111000110;     //287pi/512
   m_sin[288]  =  14'b11000000000001;     //288pi/512
   m_cos[288]  =  14'b11111110110000;     //288pi/512
   m_sin[289]  =  14'b11000000000001;     //289pi/512
   m_cos[289]  =  14'b11111110011001;     //289pi/512
   m_sin[290]  =  14'b11000000000010;     //290pi/512
   m_cos[290]  =  14'b11111110000010;     //290pi/512
   m_sin[291]  =  14'b11000000000011;     //291pi/512
   m_cos[291]  =  14'b11111101101100;     //291pi/512
   m_sin[292]  =  14'b11000000000100;     //292pi/512
   m_cos[292]  =  14'b11111101010101;     //292pi/512
   m_sin[293]  =  14'b11000000000101;     //293pi/512
   m_cos[293]  =  14'b11111100111111;     //293pi/512
   m_sin[294]  =  14'b11000000000110;     //294pi/512
   m_cos[294]  =  14'b11111100101000;     //294pi/512
   m_sin[295]  =  14'b11000000000111;     //295pi/512
   m_cos[295]  =  14'b11111100010001;     //295pi/512
   m_sin[296]  =  14'b11000000001000;     //296pi/512
   m_cos[296]  =  14'b11111011111011;     //296pi/512
   m_sin[297]  =  14'b11000000001010;     //297pi/512
   m_cos[297]  =  14'b11111011100100;     //297pi/512
   m_sin[298]  =  14'b11000000001011;     //298pi/512
   m_cos[298]  =  14'b11111011001110;     //298pi/512
   m_sin[299]  =  14'b11000000001101;     //299pi/512
   m_cos[299]  =  14'b11111010110111;     //299pi/512
   m_sin[300]  =  14'b11000000001111;     //300pi/512
   m_cos[300]  =  14'b11111010100001;     //300pi/512
   m_sin[301]  =  14'b11000000010001;     //301pi/512
   m_cos[301]  =  14'b11111010001010;     //301pi/512
   m_sin[302]  =  14'b11000000010011;     //302pi/512
   m_cos[302]  =  14'b11111001110100;     //302pi/512
   m_sin[303]  =  14'b11000000010101;     //303pi/512
   m_cos[303]  =  14'b11111001011101;     //303pi/512
   m_sin[304]  =  14'b11000000011000;     //304pi/512
   m_cos[304]  =  14'b11111001000111;     //304pi/512
   m_sin[305]  =  14'b11000000011010;     //305pi/512
   m_cos[305]  =  14'b11111000110000;     //305pi/512
   m_sin[306]  =  14'b11000000011101;     //306pi/512
   m_cos[306]  =  14'b11111000011010;     //306pi/512
   m_sin[307]  =  14'b11000000100000;     //307pi/512
   m_cos[307]  =  14'b11111000000011;     //307pi/512
   m_sin[308]  =  14'b11000000100011;     //308pi/512
   m_cos[308]  =  14'b11110111101101;     //308pi/512
   m_sin[309]  =  14'b11000000100110;     //309pi/512
   m_cos[309]  =  14'b11110111010110;     //309pi/512
   m_sin[310]  =  14'b11000000101001;     //310pi/512
   m_cos[310]  =  14'b11110111000000;     //310pi/512
   m_sin[311]  =  14'b11000000101100;     //311pi/512
   m_cos[311]  =  14'b11110110101001;     //311pi/512
   m_sin[312]  =  14'b11000000101111;     //312pi/512
   m_cos[312]  =  14'b11110110010011;     //312pi/512
   m_sin[313]  =  14'b11000000110011;     //313pi/512
   m_cos[313]  =  14'b11110101111101;     //313pi/512
   m_sin[314]  =  14'b11000000110110;     //314pi/512
   m_cos[314]  =  14'b11110101100110;     //314pi/512
   m_sin[315]  =  14'b11000000111010;     //315pi/512
   m_cos[315]  =  14'b11110101010000;     //315pi/512
   m_sin[316]  =  14'b11000000111110;     //316pi/512
   m_cos[316]  =  14'b11110100111010;     //316pi/512
   m_sin[317]  =  14'b11000001000010;     //317pi/512
   m_cos[317]  =  14'b11110100100100;     //317pi/512
   m_sin[318]  =  14'b11000001000110;     //318pi/512
   m_cos[318]  =  14'b11110100001101;     //318pi/512
   m_sin[319]  =  14'b11000001001010;     //319pi/512
   m_cos[319]  =  14'b11110011110111;     //319pi/512
   m_sin[320]  =  14'b11000001001111;     //320pi/512
   m_cos[320]  =  14'b11110011100001;     //320pi/512
   m_sin[321]  =  14'b11000001010011;     //321pi/512
   m_cos[321]  =  14'b11110011001011;     //321pi/512
   m_sin[322]  =  14'b11000001011000;     //322pi/512
   m_cos[322]  =  14'b11110010110101;     //322pi/512
   m_sin[323]  =  14'b11000001011100;     //323pi/512
   m_cos[323]  =  14'b11110010011110;     //323pi/512
   m_sin[324]  =  14'b11000001100001;     //324pi/512
   m_cos[324]  =  14'b11110010001000;     //324pi/512
   m_sin[325]  =  14'b11000001100110;     //325pi/512
   m_cos[325]  =  14'b11110001110010;     //325pi/512
   m_sin[326]  =  14'b11000001101011;     //326pi/512
   m_cos[326]  =  14'b11110001011100;     //326pi/512
   m_sin[327]  =  14'b11000001110001;     //327pi/512
   m_cos[327]  =  14'b11110001000110;     //327pi/512
   m_sin[328]  =  14'b11000001110110;     //328pi/512
   m_cos[328]  =  14'b11110000110000;     //328pi/512
   m_sin[329]  =  14'b11000001111011;     //329pi/512
   m_cos[329]  =  14'b11110000011010;     //329pi/512
   m_sin[330]  =  14'b11000010000001;     //330pi/512
   m_cos[330]  =  14'b11110000000100;     //330pi/512
   m_sin[331]  =  14'b11000010000111;     //331pi/512
   m_cos[331]  =  14'b11101111101111;     //331pi/512
   m_sin[332]  =  14'b11000010001100;     //332pi/512
   m_cos[332]  =  14'b11101111011001;     //332pi/512
   m_sin[333]  =  14'b11000010010010;     //333pi/512
   m_cos[333]  =  14'b11101111000011;     //333pi/512
   m_sin[334]  =  14'b11000010011000;     //334pi/512
   m_cos[334]  =  14'b11101110101101;     //334pi/512
   m_sin[335]  =  14'b11000010011111;     //335pi/512
   m_cos[335]  =  14'b11101110010111;     //335pi/512
   m_sin[336]  =  14'b11000010100101;     //336pi/512
   m_cos[336]  =  14'b11101110000010;     //336pi/512
   m_sin[337]  =  14'b11000010101011;     //337pi/512
   m_cos[337]  =  14'b11101101101100;     //337pi/512
   m_sin[338]  =  14'b11000010110010;     //338pi/512
   m_cos[338]  =  14'b11101101010110;     //338pi/512
   m_sin[339]  =  14'b11000010111000;     //339pi/512
   m_cos[339]  =  14'b11101101000001;     //339pi/512
   m_sin[340]  =  14'b11000010111111;     //340pi/512
   m_cos[340]  =  14'b11101100101011;     //340pi/512
   m_sin[341]  =  14'b11000011000110;     //341pi/512
   m_cos[341]  =  14'b11101100010101;     //341pi/512
   m_sin[342]  =  14'b11000011001101;     //342pi/512
   m_cos[342]  =  14'b11101100000000;     //342pi/512
   m_sin[343]  =  14'b11000011010100;     //343pi/512
   m_cos[343]  =  14'b11101011101010;     //343pi/512
   m_sin[344]  =  14'b11000011011100;     //344pi/512
   m_cos[344]  =  14'b11101011010101;     //344pi/512
   m_sin[345]  =  14'b11000011100011;     //345pi/512
   m_cos[345]  =  14'b11101011000000;     //345pi/512
   m_sin[346]  =  14'b11000011101010;     //346pi/512
   m_cos[346]  =  14'b11101010101010;     //346pi/512
   m_sin[347]  =  14'b11000011110010;     //347pi/512
   m_cos[347]  =  14'b11101010010101;     //347pi/512
   m_sin[348]  =  14'b11000011111010;     //348pi/512
   m_cos[348]  =  14'b11101010000000;     //348pi/512
   m_sin[349]  =  14'b11000100000010;     //349pi/512
   m_cos[349]  =  14'b11101001101011;     //349pi/512
   m_sin[350]  =  14'b11000100001001;     //350pi/512
   m_cos[350]  =  14'b11101001010101;     //350pi/512
   m_sin[351]  =  14'b11000100010010;     //351pi/512
   m_cos[351]  =  14'b11101001000000;     //351pi/512
   m_sin[352]  =  14'b11000100011010;     //352pi/512
   m_cos[352]  =  14'b11101000101011;     //352pi/512
   m_sin[353]  =  14'b11000100100010;     //353pi/512
   m_cos[353]  =  14'b11101000010110;     //353pi/512
   m_sin[354]  =  14'b11000100101010;     //354pi/512
   m_cos[354]  =  14'b11101000000001;     //354pi/512
   m_sin[355]  =  14'b11000100110011;     //355pi/512
   m_cos[355]  =  14'b11100111101100;     //355pi/512
   m_sin[356]  =  14'b11000100111100;     //356pi/512
   m_cos[356]  =  14'b11100111010111;     //356pi/512
   m_sin[357]  =  14'b11000101000100;     //357pi/512
   m_cos[357]  =  14'b11100111000010;     //357pi/512
   m_sin[358]  =  14'b11000101001101;     //358pi/512
   m_cos[358]  =  14'b11100110101110;     //358pi/512
   m_sin[359]  =  14'b11000101010110;     //359pi/512
   m_cos[359]  =  14'b11100110011001;     //359pi/512
   m_sin[360]  =  14'b11000101011111;     //360pi/512
   m_cos[360]  =  14'b11100110000100;     //360pi/512
   m_sin[361]  =  14'b11000101101001;     //361pi/512
   m_cos[361]  =  14'b11100101101111;     //361pi/512
   m_sin[362]  =  14'b11000101110010;     //362pi/512
   m_cos[362]  =  14'b11100101011011;     //362pi/512
   m_sin[363]  =  14'b11000101111011;     //363pi/512
   m_cos[363]  =  14'b11100101000110;     //363pi/512
   m_sin[364]  =  14'b11000110000101;     //364pi/512
   m_cos[364]  =  14'b11100100110010;     //364pi/512
   m_sin[365]  =  14'b11000110001111;     //365pi/512
   m_cos[365]  =  14'b11100100011101;     //365pi/512
   m_sin[366]  =  14'b11000110011000;     //366pi/512
   m_cos[366]  =  14'b11100100001001;     //366pi/512
   m_sin[367]  =  14'b11000110100010;     //367pi/512
   m_cos[367]  =  14'b11100011110101;     //367pi/512
   m_sin[368]  =  14'b11000110101100;     //368pi/512
   m_cos[368]  =  14'b11100011100000;     //368pi/512
   m_sin[369]  =  14'b11000110110110;     //369pi/512
   m_cos[369]  =  14'b11100011001100;     //369pi/512
   m_sin[370]  =  14'b11000111000001;     //370pi/512
   m_cos[370]  =  14'b11100010111000;     //370pi/512
   m_sin[371]  =  14'b11000111001011;     //371pi/512
   m_cos[371]  =  14'b11100010100100;     //371pi/512
   m_sin[372]  =  14'b11000111010110;     //372pi/512
   m_cos[372]  =  14'b11100010010000;     //372pi/512
   m_sin[373]  =  14'b11000111100000;     //373pi/512
   m_cos[373]  =  14'b11100001111100;     //373pi/512
   m_sin[374]  =  14'b11000111101011;     //374pi/512
   m_cos[374]  =  14'b11100001101000;     //374pi/512
   m_sin[375]  =  14'b11000111110110;     //375pi/512
   m_cos[375]  =  14'b11100001010100;     //375pi/512
   m_sin[376]  =  14'b11001000000000;     //376pi/512
   m_cos[376]  =  14'b11100001000000;     //376pi/512
   m_sin[377]  =  14'b11001000001011;     //377pi/512
   m_cos[377]  =  14'b11100000101100;     //377pi/512
   m_sin[378]  =  14'b11001000010111;     //378pi/512
   m_cos[378]  =  14'b11100000011001;     //378pi/512
   m_sin[379]  =  14'b11001000100010;     //379pi/512
   m_cos[379]  =  14'b11100000000101;     //379pi/512
   m_sin[380]  =  14'b11001000101101;     //380pi/512
   m_cos[380]  =  14'b11011111110010;     //380pi/512
   m_sin[381]  =  14'b11001000111001;     //381pi/512
   m_cos[381]  =  14'b11011111011110;     //381pi/512
   m_sin[382]  =  14'b11001001000100;     //382pi/512
   m_cos[382]  =  14'b11011111001011;     //382pi/512
   m_sin[383]  =  14'b11001001010000;     //383pi/512
   m_cos[383]  =  14'b11011110110111;     //383pi/512
   m_sin[384]  =  14'b11001001011100;     //384pi/512
   m_cos[384]  =  14'b11011110100100;     //384pi/512
   m_sin[385]  =  14'b11001001100111;     //385pi/512
   m_cos[385]  =  14'b11011110010001;     //385pi/512
   m_sin[386]  =  14'b11001001110011;     //386pi/512
   m_cos[386]  =  14'b11011101111101;     //386pi/512
   m_sin[387]  =  14'b11001010000000;     //387pi/512
   m_cos[387]  =  14'b11011101101010;     //387pi/512
   m_sin[388]  =  14'b11001010001100;     //388pi/512
   m_cos[388]  =  14'b11011101010111;     //388pi/512
   m_sin[389]  =  14'b11001010011000;     //389pi/512
   m_cos[389]  =  14'b11011101000100;     //389pi/512
   m_sin[390]  =  14'b11001010100100;     //390pi/512
   m_cos[390]  =  14'b11011100110001;     //390pi/512
   m_sin[391]  =  14'b11001010110001;     //391pi/512
   m_cos[391]  =  14'b11011100011110;     //391pi/512
   m_sin[392]  =  14'b11001010111110;     //392pi/512
   m_cos[392]  =  14'b11011100001100;     //392pi/512
   m_sin[393]  =  14'b11001011001010;     //393pi/512
   m_cos[393]  =  14'b11011011111001;     //393pi/512
   m_sin[394]  =  14'b11001011010111;     //394pi/512
   m_cos[394]  =  14'b11011011100110;     //394pi/512
   m_sin[395]  =  14'b11001011100100;     //395pi/512
   m_cos[395]  =  14'b11011011010100;     //395pi/512
   m_sin[396]  =  14'b11001011110001;     //396pi/512
   m_cos[396]  =  14'b11011011000001;     //396pi/512
   m_sin[397]  =  14'b11001011111110;     //397pi/512
   m_cos[397]  =  14'b11011010101111;     //397pi/512
   m_sin[398]  =  14'b11001100001011;     //398pi/512
   m_cos[398]  =  14'b11011010011100;     //398pi/512
   m_sin[399]  =  14'b11001100011001;     //399pi/512
   m_cos[399]  =  14'b11011010001010;     //399pi/512
   m_sin[400]  =  14'b11001100100110;     //400pi/512
   m_cos[400]  =  14'b11011001111000;     //400pi/512
   m_sin[401]  =  14'b11001100110100;     //401pi/512
   m_cos[401]  =  14'b11011001100110;     //401pi/512
   m_sin[402]  =  14'b11001101000001;     //402pi/512
   m_cos[402]  =  14'b11011001010100;     //402pi/512
   m_sin[403]  =  14'b11001101001111;     //403pi/512
   m_cos[403]  =  14'b11011001000010;     //403pi/512
   m_sin[404]  =  14'b11001101011101;     //404pi/512
   m_cos[404]  =  14'b11011000110000;     //404pi/512
   m_sin[405]  =  14'b11001101101011;     //405pi/512
   m_cos[405]  =  14'b11011000011110;     //405pi/512
   m_sin[406]  =  14'b11001101111001;     //406pi/512
   m_cos[406]  =  14'b11011000001100;     //406pi/512
   m_sin[407]  =  14'b11001110000111;     //407pi/512
   m_cos[407]  =  14'b11010111111011;     //407pi/512
   m_sin[408]  =  14'b11001110010101;     //408pi/512
   m_cos[408]  =  14'b11010111101001;     //408pi/512
   m_sin[409]  =  14'b11001110100011;     //409pi/512
   m_cos[409]  =  14'b11010111011000;     //409pi/512
   m_sin[410]  =  14'b11001110110010;     //410pi/512
   m_cos[410]  =  14'b11010111000110;     //410pi/512
   m_sin[411]  =  14'b11001111000000;     //411pi/512
   m_cos[411]  =  14'b11010110110101;     //411pi/512
   m_sin[412]  =  14'b11001111001111;     //412pi/512
   m_cos[412]  =  14'b11010110100100;     //412pi/512
   m_sin[413]  =  14'b11001111011110;     //413pi/512
   m_cos[413]  =  14'b11010110010010;     //413pi/512
   m_sin[414]  =  14'b11001111101100;     //414pi/512
   m_cos[414]  =  14'b11010110000001;     //414pi/512
   m_sin[415]  =  14'b11001111111011;     //415pi/512
   m_cos[415]  =  14'b11010101110000;     //415pi/512
   m_sin[416]  =  14'b11010000001010;     //416pi/512
   m_cos[416]  =  14'b11010101011111;     //416pi/512
   m_sin[417]  =  14'b11010000011001;     //417pi/512
   m_cos[417]  =  14'b11010101001110;     //417pi/512
   m_sin[418]  =  14'b11010000101000;     //418pi/512
   m_cos[418]  =  14'b11010100111110;     //418pi/512
   m_sin[419]  =  14'b11010000111000;     //419pi/512
   m_cos[419]  =  14'b11010100101101;     //419pi/512
   m_sin[420]  =  14'b11010001000111;     //420pi/512
   m_cos[420]  =  14'b11010100011100;     //420pi/512
   m_sin[421]  =  14'b11010001010110;     //421pi/512
   m_cos[421]  =  14'b11010100001100;     //421pi/512
   m_sin[422]  =  14'b11010001100110;     //422pi/512
   m_cos[422]  =  14'b11010011111011;     //422pi/512
   m_sin[423]  =  14'b11010001110110;     //423pi/512
   m_cos[423]  =  14'b11010011101011;     //423pi/512
   m_sin[424]  =  14'b11010010000101;     //424pi/512
   m_cos[424]  =  14'b11010011011011;     //424pi/512
   m_sin[425]  =  14'b11010010010101;     //425pi/512
   m_cos[425]  =  14'b11010011001010;     //425pi/512
   m_sin[426]  =  14'b11010010100101;     //426pi/512
   m_cos[426]  =  14'b11010010111010;     //426pi/512
   m_sin[427]  =  14'b11010010110101;     //427pi/512
   m_cos[427]  =  14'b11010010101010;     //427pi/512
   m_sin[428]  =  14'b11010011000101;     //428pi/512
   m_cos[428]  =  14'b11010010011010;     //428pi/512
   m_sin[429]  =  14'b11010011010101;     //429pi/512
   m_cos[429]  =  14'b11010010001011;     //429pi/512
   m_sin[430]  =  14'b11010011100101;     //430pi/512
   m_cos[430]  =  14'b11010001111011;     //430pi/512
   m_sin[431]  =  14'b11010011110110;     //431pi/512
   m_cos[431]  =  14'b11010001101011;     //431pi/512
   m_sin[432]  =  14'b11010100000110;     //432pi/512
   m_cos[432]  =  14'b11010001011100;     //432pi/512
   m_sin[433]  =  14'b11010100010111;     //433pi/512
   m_cos[433]  =  14'b11010001001100;     //433pi/512
   m_sin[434]  =  14'b11010100100111;     //434pi/512
   m_cos[434]  =  14'b11010000111101;     //434pi/512
   m_sin[435]  =  14'b11010100111000;     //435pi/512
   m_cos[435]  =  14'b11010000101110;     //435pi/512
   m_sin[436]  =  14'b11010101001001;     //436pi/512
   m_cos[436]  =  14'b11010000011110;     //436pi/512
   m_sin[437]  =  14'b11010101011010;     //437pi/512
   m_cos[437]  =  14'b11010000001111;     //437pi/512
   m_sin[438]  =  14'b11010101101011;     //438pi/512
   m_cos[438]  =  14'b11010000000000;     //438pi/512
   m_sin[439]  =  14'b11010101111100;     //439pi/512
   m_cos[439]  =  14'b11001111110001;     //439pi/512
   m_sin[440]  =  14'b11010110001101;     //440pi/512
   m_cos[440]  =  14'b11001111100010;     //440pi/512
   m_sin[441]  =  14'b11010110011110;     //441pi/512
   m_cos[441]  =  14'b11001111010100;     //441pi/512
   m_sin[442]  =  14'b11010110101111;     //442pi/512
   m_cos[442]  =  14'b11001111000101;     //442pi/512
   m_sin[443]  =  14'b11010111000000;     //443pi/512
   m_cos[443]  =  14'b11001110110111;     //443pi/512
   m_sin[444]  =  14'b11010111010010;     //444pi/512
   m_cos[444]  =  14'b11001110101000;     //444pi/512
   m_sin[445]  =  14'b11010111100011;     //445pi/512
   m_cos[445]  =  14'b11001110011010;     //445pi/512
   m_sin[446]  =  14'b11010111110101;     //446pi/512
   m_cos[446]  =  14'b11001110001100;     //446pi/512
   m_sin[447]  =  14'b11011000000110;     //447pi/512
   m_cos[447]  =  14'b11001101111101;     //447pi/512
   m_sin[448]  =  14'b11011000011000;     //448pi/512
   m_cos[448]  =  14'b11001101101111;     //448pi/512
   m_sin[449]  =  14'b11011000101010;     //449pi/512
   m_cos[449]  =  14'b11001101100001;     //449pi/512
   m_sin[450]  =  14'b11011000111100;     //450pi/512
   m_cos[450]  =  14'b11001101010100;     //450pi/512
   m_sin[451]  =  14'b11011001001110;     //451pi/512
   m_cos[451]  =  14'b11001101000110;     //451pi/512
   m_sin[452]  =  14'b11011001100000;     //452pi/512
   m_cos[452]  =  14'b11001100111000;     //452pi/512
   m_sin[453]  =  14'b11011001110010;     //453pi/512
   m_cos[453]  =  14'b11001100101011;     //453pi/512
   m_sin[454]  =  14'b11011010000100;     //454pi/512
   m_cos[454]  =  14'b11001100011101;     //454pi/512
   m_sin[455]  =  14'b11011010010110;     //455pi/512
   m_cos[455]  =  14'b11001100010000;     //455pi/512
   m_sin[456]  =  14'b11011010101001;     //456pi/512
   m_cos[456]  =  14'b11001100000010;     //456pi/512
   m_sin[457]  =  14'b11011010111011;     //457pi/512
   m_cos[457]  =  14'b11001011110101;     //457pi/512
   m_sin[458]  =  14'b11011011001110;     //458pi/512
   m_cos[458]  =  14'b11001011101000;     //458pi/512
   m_sin[459]  =  14'b11011011100000;     //459pi/512
   m_cos[459]  =  14'b11001011011011;     //459pi/512
   m_sin[460]  =  14'b11011011110011;     //460pi/512
   m_cos[460]  =  14'b11001011001110;     //460pi/512
   m_sin[461]  =  14'b11011100000101;     //461pi/512
   m_cos[461]  =  14'b11001011000010;     //461pi/512
   m_sin[462]  =  14'b11011100011000;     //462pi/512
   m_cos[462]  =  14'b11001010110101;     //462pi/512
   m_sin[463]  =  14'b11011100101011;     //463pi/512
   m_cos[463]  =  14'b11001010101001;     //463pi/512
   m_sin[464]  =  14'b11011100111110;     //464pi/512
   m_cos[464]  =  14'b11001010011100;     //464pi/512
   m_sin[465]  =  14'b11011101010001;     //465pi/512
   m_cos[465]  =  14'b11001010010000;     //465pi/512
   m_sin[466]  =  14'b11011101100100;     //466pi/512
   m_cos[466]  =  14'b11001010000100;     //466pi/512
   m_sin[467]  =  14'b11011101110111;     //467pi/512
   m_cos[467]  =  14'b11001001110111;     //467pi/512
   m_sin[468]  =  14'b11011110001010;     //468pi/512
   m_cos[468]  =  14'b11001001101011;     //468pi/512
   m_sin[469]  =  14'b11011110011101;     //469pi/512
   m_cos[469]  =  14'b11001001100000;     //469pi/512
   m_sin[470]  =  14'b11011110110001;     //470pi/512
   m_cos[470]  =  14'b11001001010100;     //470pi/512
   m_sin[471]  =  14'b11011111000100;     //471pi/512
   m_cos[471]  =  14'b11001001001000;     //471pi/512
   m_sin[472]  =  14'b11011111011000;     //472pi/512
   m_cos[472]  =  14'b11001000111100;     //472pi/512
   m_sin[473]  =  14'b11011111101011;     //473pi/512
   m_cos[473]  =  14'b11001000110001;     //473pi/512
   m_sin[474]  =  14'b11011111111111;     //474pi/512
   m_cos[474]  =  14'b11001000100110;     //474pi/512
   m_sin[475]  =  14'b11100000010010;     //475pi/512
   m_cos[475]  =  14'b11001000011010;     //475pi/512
   m_sin[476]  =  14'b11100000100110;     //476pi/512
   m_cos[476]  =  14'b11001000001111;     //476pi/512
   m_sin[477]  =  14'b11100000111010;     //477pi/512
   m_cos[477]  =  14'b11001000000100;     //477pi/512
   m_sin[478]  =  14'b11100001001101;     //478pi/512
   m_cos[478]  =  14'b11000111111001;     //478pi/512
   m_sin[479]  =  14'b11100001100001;     //479pi/512
   m_cos[479]  =  14'b11000111101110;     //479pi/512
   m_sin[480]  =  14'b11100001110101;     //480pi/512
   m_cos[480]  =  14'b11000111100100;     //480pi/512
   m_sin[481]  =  14'b11100010001001;     //481pi/512
   m_cos[481]  =  14'b11000111011001;     //481pi/512
   m_sin[482]  =  14'b11100010011101;     //482pi/512
   m_cos[482]  =  14'b11000111001111;     //482pi/512
   m_sin[483]  =  14'b11100010110001;     //483pi/512
   m_cos[483]  =  14'b11000111000100;     //483pi/512
   m_sin[484]  =  14'b11100011000101;     //484pi/512
   m_cos[484]  =  14'b11000110111010;     //484pi/512
   m_sin[485]  =  14'b11100011011010;     //485pi/512
   m_cos[485]  =  14'b11000110110000;     //485pi/512
   m_sin[486]  =  14'b11100011101110;     //486pi/512
   m_cos[486]  =  14'b11000110100110;     //486pi/512
   m_sin[487]  =  14'b11100100000010;     //487pi/512
   m_cos[487]  =  14'b11000110011100;     //487pi/512
   m_sin[488]  =  14'b11100100010111;     //488pi/512
   m_cos[488]  =  14'b11000110010010;     //488pi/512
   m_sin[489]  =  14'b11100100101011;     //489pi/512
   m_cos[489]  =  14'b11000110001000;     //489pi/512
   m_sin[490]  =  14'b11100100111111;     //490pi/512
   m_cos[490]  =  14'b11000101111111;     //490pi/512
   m_sin[491]  =  14'b11100101010100;     //491pi/512
   m_cos[491]  =  14'b11000101110101;     //491pi/512
   m_sin[492]  =  14'b11100101101001;     //492pi/512
   m_cos[492]  =  14'b11000101101100;     //492pi/512
   m_sin[493]  =  14'b11100101111101;     //493pi/512
   m_cos[493]  =  14'b11000101100010;     //493pi/512
   m_sin[494]  =  14'b11100110010010;     //494pi/512
   m_cos[494]  =  14'b11000101011001;     //494pi/512
   m_sin[495]  =  14'b11100110100111;     //495pi/512
   m_cos[495]  =  14'b11000101010000;     //495pi/512
   m_sin[496]  =  14'b11100110111011;     //496pi/512
   m_cos[496]  =  14'b11000101000111;     //496pi/512
   m_sin[497]  =  14'b11100111010000;     //497pi/512
   m_cos[497]  =  14'b11000100111111;     //497pi/512
   m_sin[498]  =  14'b11100111100101;     //498pi/512
   m_cos[498]  =  14'b11000100110110;     //498pi/512
   m_sin[499]  =  14'b11100111111010;     //499pi/512
   m_cos[499]  =  14'b11000100101101;     //499pi/512
   m_sin[500]  =  14'b11101000001111;     //500pi/512
   m_cos[500]  =  14'b11000100100101;     //500pi/512
   m_sin[501]  =  14'b11101000100100;     //501pi/512
   m_cos[501]  =  14'b11000100011100;     //501pi/512
   m_sin[502]  =  14'b11101000111001;     //502pi/512
   m_cos[502]  =  14'b11000100010100;     //502pi/512
   m_sin[503]  =  14'b11101001001110;     //503pi/512
   m_cos[503]  =  14'b11000100001100;     //503pi/512
   m_sin[504]  =  14'b11101001100011;     //504pi/512
   m_cos[504]  =  14'b11000100000100;     //504pi/512
   m_sin[505]  =  14'b11101001111001;     //505pi/512
   m_cos[505]  =  14'b11000011111100;     //505pi/512
   m_sin[506]  =  14'b11101010001110;     //506pi/512
   m_cos[506]  =  14'b11000011110101;     //506pi/512
   m_sin[507]  =  14'b11101010100011;     //507pi/512
   m_cos[507]  =  14'b11000011101101;     //507pi/512
   m_sin[508]  =  14'b11101010111001;     //508pi/512
   m_cos[508]  =  14'b11000011100101;     //508pi/512
   m_sin[509]  =  14'b11101011001110;     //509pi/512
   m_cos[509]  =  14'b11000011011110;     //509pi/512
   m_sin[510]  =  14'b11101011100011;     //510pi/512
   m_cos[510]  =  14'b11000011010111;     //510pi/512
   m_sin[511]  =  14'b11101011111001;     //511pi/512
   m_cos[511]  =  14'b11000011010000;     //511pi/512
end

endmodule