module  M_TWIDLE_16_bit #(parameter SIZE =10, word_length_tw = 16) (
    input            clk,
    input            en_rd, 
    input   [10:0]   rd_ptr_angle,
    input            en_modf, 

    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );


reg signed [word_length_tw-1:0]  cos  [511:0];
reg signed [word_length_tw-1:0]  sin  [511:0];

reg signed [word_length_tw-1:0]  m_cos  [511:0];
reg signed [word_length_tw-1:0]  m_sin  [511:0];

reg signed [word_length_tw-1:0]  cos_temp;
reg signed [word_length_tw-1:0]  sin_temp;

reg signed [word_length_tw-1:0]  m_cos_temp;
reg signed [word_length_tw-1:0]  m_sin_temp;


//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & ~ en_modf ) begin
                  cos_temp           <= cos   [rd_ptr_angle];
                  sin_temp           <= sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & en_modf ) begin
                  m_cos_temp           <= m_cos   [rd_ptr_angle];
                  m_sin_temp           <= m_sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(*) begin 
             if (en_modf ) begin
                  cos_data           <= m_cos_temp;
                  sin_data           <= m_sin_temp;
             end else begin
                  cos_data           <= cos_temp;
                  sin_data           <= sin_temp;
             end
        end
//----------------------------------------------------------------------------------------
initial begin
   sin[0]  =  16'b0000_0000_0000_0000;     //0pi/512
   cos[0]  =  16'b0100_0000_0000_0000;     //0pi/512
   sin[1]  =  16'b1111_1111_1001_1011;     //1pi/512
   cos[1]  =  16'b0011_1111_1111_1111;     //1pi/512
   sin[2]  =  16'b1111_1111_0011_0111;     //2pi/512
   cos[2]  =  16'b0011_1111_1111_1110;     //2pi/512
   sin[3]  =  16'b1111_1110_1101_0010;     //3pi/512
   cos[3]  =  16'b0011_1111_1111_1101;     //3pi/512
   sin[4]  =  16'b1111_1110_0110_1110;     //4pi/512
   cos[4]  =  16'b0011_1111_1111_1011;     //4pi/512
   sin[5]  =  16'b1111_1110_0000_1001;     //5pi/512
   cos[5]  =  16'b0011_1111_1111_1000;     //5pi/512
   sin[6]  =  16'b1111_1101_1010_0101;     //6pi/512
   cos[6]  =  16'b0011_1111_1111_0100;     //6pi/512
   sin[7]  =  16'b1111_1101_0100_0000;     //7pi/512
   cos[7]  =  16'b0011_1111_1111_0000;     //7pi/512
   sin[8]  =  16'b1111_1100_1101_1100;     //8pi/512
   cos[8]  =  16'b0011_1111_1110_1100;     //8pi/512
   sin[9]  =  16'b1111_1100_0111_1000;     //9pi/512
   cos[9]  =  16'b0011_1111_1110_0111;     //9pi/512
   sin[10]  =  16'b1111_1100_0001_0011;     //10pi/512
   cos[10]  =  16'b0011_1111_1110_0001;     //10pi/512
   sin[11]  =  16'b1111_1011_1010_1111;     //11pi/512
   cos[11]  =  16'b0011_1111_1101_1010;     //11pi/512
   sin[12]  =  16'b1111_1011_0100_1011;     //12pi/512
   cos[12]  =  16'b0011_1111_1101_0011;     //12pi/512
   sin[13]  =  16'b1111_1010_1110_0110;     //13pi/512
   cos[13]  =  16'b0011_1111_1100_1011;     //13pi/512
   sin[14]  =  16'b1111_1010_1000_0010;     //14pi/512
   cos[14]  =  16'b0011_1111_1100_0011;     //14pi/512
   sin[15]  =  16'b1111_1010_0001_1110;     //15pi/512
   cos[15]  =  16'b0011_1111_1011_1010;     //15pi/512
   sin[16]  =  16'b1111_1001_1011_1010;     //16pi/512
   cos[16]  =  16'b0011_1111_1011_0001;     //16pi/512
   sin[17]  =  16'b1111_1001_0101_0110;     //17pi/512
   cos[17]  =  16'b0011_1111_1010_0110;     //17pi/512
   sin[18]  =  16'b1111_1000_1111_0010;     //18pi/512
   cos[18]  =  16'b0011_1111_1001_1100;     //18pi/512
   sin[19]  =  16'b1111_1000_1000_1110;     //19pi/512
   cos[19]  =  16'b0011_1111_1001_0000;     //19pi/512
   sin[20]  =  16'b1111_1000_0010_1010;     //20pi/512
   cos[20]  =  16'b0011_1111_1000_0100;     //20pi/512
   sin[21]  =  16'b1111_0111_1100_0111;     //21pi/512
   cos[21]  =  16'b0011_1111_0111_1000;     //21pi/512
   sin[22]  =  16'b1111_0111_0110_0011;     //22pi/512
   cos[22]  =  16'b0011_1111_0110_1010;     //22pi/512
   sin[23]  =  16'b1111_0110_1111_1111;     //23pi/512
   cos[23]  =  16'b0011_1111_0101_1101;     //23pi/512
   sin[24]  =  16'b1111_0110_1001_1100;     //24pi/512
   cos[24]  =  16'b0011_1111_0100_1110;     //24pi/512
   sin[25]  =  16'b1111_0110_0011_1001;     //25pi/512
   cos[25]  =  16'b0011_1111_0011_1111;     //25pi/512
   sin[26]  =  16'b1111_0101_1101_0101;     //26pi/512
   cos[26]  =  16'b0011_1111_0010_1111;     //26pi/512
   sin[27]  =  16'b1111_0101_0111_0010;     //27pi/512
   cos[27]  =  16'b0011_1111_0001_1111;     //27pi/512
   sin[28]  =  16'b1111_0101_0000_1111;     //28pi/512
   cos[28]  =  16'b0011_1111_0000_1110;     //28pi/512
   sin[29]  =  16'b1111_0100_1010_1100;     //29pi/512
   cos[29]  =  16'b0011_1110_1111_1101;     //29pi/512
   sin[30]  =  16'b1111_0100_0100_1001;     //30pi/512
   cos[30]  =  16'b0011_1110_1110_1011;     //30pi/512
   sin[31]  =  16'b1111_0011_1110_0110;     //31pi/512
   cos[31]  =  16'b0011_1110_1101_1000;     //31pi/512
   sin[32]  =  16'b1111_0011_1000_0100;     //32pi/512
   cos[32]  =  16'b0011_1110_1100_0101;     //32pi/512
   sin[33]  =  16'b1111_0011_0010_0001;     //33pi/512
   cos[33]  =  16'b0011_1110_1011_0001;     //33pi/512
   sin[34]  =  16'b1111_0010_1011_1111;     //34pi/512
   cos[34]  =  16'b0011_1110_1001_1100;     //34pi/512
   sin[35]  =  16'b1111_0010_0101_1100;     //35pi/512
   cos[35]  =  16'b0011_1110_1000_0111;     //35pi/512
   sin[36]  =  16'b1111_0001_1111_1010;     //36pi/512
   cos[36]  =  16'b0011_1110_0111_0001;     //36pi/512
   sin[37]  =  16'b1111_0001_1001_1000;     //37pi/512
   cos[37]  =  16'b0011_1110_0101_1011;     //37pi/512
   sin[38]  =  16'b1111_0001_0011_0110;     //38pi/512
   cos[38]  =  16'b0011_1110_0100_0100;     //38pi/512
   sin[39]  =  16'b1111_0000_1101_0101;     //39pi/512
   cos[39]  =  16'b0011_1110_0010_1101;     //39pi/512
   sin[40]  =  16'b1111_0000_0111_0011;     //40pi/512
   cos[40]  =  16'b0011_1110_0001_0100;     //40pi/512
   sin[41]  =  16'b1111_0000_0001_0010;     //41pi/512
   cos[41]  =  16'b0011_1101_1111_1100;     //41pi/512
   sin[42]  =  16'b1110_1111_1011_0000;     //42pi/512
   cos[42]  =  16'b0011_1101_1110_0010;     //42pi/512
   sin[43]  =  16'b1110_1111_0100_1111;     //43pi/512
   cos[43]  =  16'b0011_1101_1100_1001;     //43pi/512
   sin[44]  =  16'b1110_1110_1110_1110;     //44pi/512
   cos[44]  =  16'b0011_1101_1010_1110;     //44pi/512
   sin[45]  =  16'b1110_1110_1000_1101;     //45pi/512
   cos[45]  =  16'b0011_1101_1001_0011;     //45pi/512
   sin[46]  =  16'b1110_1110_0010_1101;     //46pi/512
   cos[46]  =  16'b0011_1101_0111_0111;     //46pi/512
   sin[47]  =  16'b1110_1101_1100_1100;     //47pi/512
   cos[47]  =  16'b0011_1101_0101_1011;     //47pi/512
   sin[48]  =  16'b1110_1101_0110_1100;     //48pi/512
   cos[48]  =  16'b0011_1101_0011_1110;     //48pi/512
   sin[49]  =  16'b1110_1101_0000_1100;     //49pi/512
   cos[49]  =  16'b0011_1101_0010_0001;     //49pi/512
   sin[50]  =  16'b1110_1100_1010_1100;     //50pi/512
   cos[50]  =  16'b0011_1101_0000_0010;     //50pi/512
   sin[51]  =  16'b1110_1100_0100_1100;     //51pi/512
   cos[51]  =  16'b0011_1100_1110_0100;     //51pi/512
   sin[52]  =  16'b1110_1011_1110_1101;     //52pi/512
   cos[52]  =  16'b0011_1100_1100_0101;     //52pi/512
   sin[53]  =  16'b1110_1011_1000_1101;     //53pi/512
   cos[53]  =  16'b0011_1100_1010_0101;     //53pi/512
   sin[54]  =  16'b1110_1011_0010_1110;     //54pi/512
   cos[54]  =  16'b0011_1100_1000_0100;     //54pi/512
   sin[55]  =  16'b1110_1010_1100_1111;     //55pi/512
   cos[55]  =  16'b0011_1100_0110_0011;     //55pi/512
   sin[56]  =  16'b1110_1010_0111_0000;     //56pi/512
   cos[56]  =  16'b0011_1100_0100_0010;     //56pi/512
   sin[57]  =  16'b1110_1010_0001_0010;     //57pi/512
   cos[57]  =  16'b0011_1100_0010_0000;     //57pi/512
   sin[58]  =  16'b1110_1001_1011_0100;     //58pi/512
   cos[58]  =  16'b0011_1011_1111_1101;     //58pi/512
   sin[59]  =  16'b1110_1001_0101_0101;     //59pi/512
   cos[59]  =  16'b0011_1011_1101_1010;     //59pi/512
   sin[60]  =  16'b1110_1000_1111_0111;     //60pi/512
   cos[60]  =  16'b0011_1011_1011_0110;     //60pi/512
   sin[61]  =  16'b1110_1000_1001_1010;     //61pi/512
   cos[61]  =  16'b0011_1011_1001_0001;     //61pi/512
   sin[62]  =  16'b1110_1000_0011_1100;     //62pi/512
   cos[62]  =  16'b0011_1011_0110_1100;     //62pi/512
   sin[63]  =  16'b1110_0111_1101_1111;     //63pi/512
   cos[63]  =  16'b0011_1011_0100_0111;     //63pi/512
   sin[64]  =  16'b1110_0111_1000_0010;     //64pi/512
   cos[64]  =  16'b0011_1011_0010_0000;     //64pi/512
   sin[65]  =  16'b1110_0111_0010_0101;     //65pi/512
   cos[65]  =  16'b0011_1010_1111_1010;     //65pi/512
   sin[66]  =  16'b1110_0110_1100_1001;     //66pi/512
   cos[66]  =  16'b0011_1010_1101_0010;     //66pi/512
   sin[67]  =  16'b1110_0110_0110_1101;     //67pi/512
   cos[67]  =  16'b0011_1010_1010_1010;     //67pi/512
   sin[68]  =  16'b1110_0110_0001_0001;     //68pi/512
   cos[68]  =  16'b0011_1010_1000_0010;     //68pi/512
   sin[69]  =  16'b1110_0101_1011_0101;     //69pi/512
   cos[69]  =  16'b0011_1010_0101_1001;     //69pi/512
   sin[70]  =  16'b1110_0101_0101_1001;     //70pi/512
   cos[70]  =  16'b0011_1010_0010_1111;     //70pi/512
   sin[71]  =  16'b1110_0100_1111_1110;     //71pi/512
   cos[71]  =  16'b0011_1010_0000_0101;     //71pi/512
   sin[72]  =  16'b1110_0100_1010_0011;     //72pi/512
   cos[72]  =  16'b0011_1001_1101_1010;     //72pi/512
   sin[73]  =  16'b1110_0100_0100_1000;     //73pi/512
   cos[73]  =  16'b0011_1001_1010_1111;     //73pi/512
   sin[74]  =  16'b1110_0011_1110_1110;     //74pi/512
   cos[74]  =  16'b0011_1001_1000_0011;     //74pi/512
   sin[75]  =  16'b1110_0011_1001_0100;     //75pi/512
   cos[75]  =  16'b0011_1001_0101_0111;     //75pi/512
   sin[76]  =  16'b1110_0011_0011_1010;     //76pi/512
   cos[76]  =  16'b0011_1001_0010_1010;     //76pi/512
   sin[77]  =  16'b1110_0010_1110_0000;     //77pi/512
   cos[77]  =  16'b0011_1000_1111_1101;     //77pi/512
   sin[78]  =  16'b1110_0010_1000_0111;     //78pi/512
   cos[78]  =  16'b0011_1000_1100_1111;     //78pi/512
   sin[79]  =  16'b1110_0010_0010_1101;     //79pi/512
   cos[79]  =  16'b0011_1000_1010_0000;     //79pi/512
   sin[80]  =  16'b1110_0001_1101_0101;     //80pi/512
   cos[80]  =  16'b0011_1000_0111_0001;     //80pi/512
   sin[81]  =  16'b1110_0001_0111_1100;     //81pi/512
   cos[81]  =  16'b0011_1000_0100_0001;     //81pi/512
   sin[82]  =  16'b1110_0001_0010_0100;     //82pi/512
   cos[82]  =  16'b0011_1000_0001_0001;     //82pi/512
   sin[83]  =  16'b1110_0000_1100_1100;     //83pi/512
   cos[83]  =  16'b0011_0111_1110_0000;     //83pi/512
   sin[84]  =  16'b1110_0000_0111_0100;     //84pi/512
   cos[84]  =  16'b0011_0111_1010_1111;     //84pi/512
   sin[85]  =  16'b1110_0000_0001_1101;     //85pi/512
   cos[85]  =  16'b0011_0111_0111_1101;     //85pi/512
   sin[86]  =  16'b1101_1111_1100_0110;     //86pi/512
   cos[86]  =  16'b0011_0111_0100_1011;     //86pi/512
   sin[87]  =  16'b1101_1111_0110_1111;     //87pi/512
   cos[87]  =  16'b0011_0111_0001_1000;     //87pi/512
   sin[88]  =  16'b1101_1111_0001_1001;     //88pi/512
   cos[88]  =  16'b0011_0110_1110_0101;     //88pi/512
   sin[89]  =  16'b1101_1110_1100_0011;     //89pi/512
   cos[89]  =  16'b0011_0110_1011_0001;     //89pi/512
   sin[90]  =  16'b1101_1110_0110_1101;     //90pi/512
   cos[90]  =  16'b0011_0110_0111_1100;     //90pi/512
   sin[91]  =  16'b1101_1110_0001_1000;     //91pi/512
   cos[91]  =  16'b0011_0110_0100_0111;     //91pi/512
   sin[92]  =  16'b1101_1101_1100_0011;     //92pi/512
   cos[92]  =  16'b0011_0110_0001_0010;     //92pi/512
   sin[93]  =  16'b1101_1101_0110_1110;     //93pi/512
   cos[93]  =  16'b0011_0101_1101_1100;     //93pi/512
   sin[94]  =  16'b1101_1101_0001_1001;     //94pi/512
   cos[94]  =  16'b0011_0101_1010_0101;     //94pi/512
   sin[95]  =  16'b1101_1100_1100_0101;     //95pi/512
   cos[95]  =  16'b0011_0101_0110_1110;     //95pi/512
   sin[96]  =  16'b1101_1100_0111_0010;     //96pi/512
   cos[96]  =  16'b0011_0101_0011_0110;     //96pi/512
   sin[97]  =  16'b1101_1100_0001_1110;     //97pi/512
   cos[97]  =  16'b0011_0100_1111_1110;     //97pi/512
   sin[98]  =  16'b1101_1011_1100_1011;     //98pi/512
   cos[98]  =  16'b0011_0100_1100_0110;     //98pi/512
   sin[99]  =  16'b1101_1011_0111_1000;     //99pi/512
   cos[99]  =  16'b0011_0100_1000_1100;     //99pi/512
   sin[100]  =  16'b1101_1011_0010_0110;     //100pi/512
   cos[100]  =  16'b0011_0100_0101_0011;     //100pi/512
   sin[101]  =  16'b1101_1010_1101_0100;     //101pi/512
   cos[101]  =  16'b0011_0100_0001_1001;     //101pi/512
   sin[102]  =  16'b1101_1010_1000_0010;     //102pi/512
   cos[102]  =  16'b0011_0011_1101_1110;     //102pi/512
   sin[103]  =  16'b1101_1010_0011_0001;     //103pi/512
   cos[103]  =  16'b0011_0011_1010_0011;     //103pi/512
   sin[104]  =  16'b1101_1001_1110_0000;     //104pi/512
   cos[104]  =  16'b0011_0011_0110_0111;     //104pi/512
   sin[105]  =  16'b1101_1001_1000_1111;     //105pi/512
   cos[105]  =  16'b0011_0011_0010_1011;     //105pi/512
   sin[106]  =  16'b1101_1001_0011_1111;     //106pi/512
   cos[106]  =  16'b0011_0010_1110_1110;     //106pi/512
   sin[107]  =  16'b1101_1000_1110_1111;     //107pi/512
   cos[107]  =  16'b0011_0010_1011_0001;     //107pi/512
   sin[108]  =  16'b1101_1000_1010_0000;     //108pi/512
   cos[108]  =  16'b0011_0010_0111_0100;     //108pi/512
   sin[109]  =  16'b1101_1000_0101_0001;     //109pi/512
   cos[109]  =  16'b0011_0010_0011_0110;     //109pi/512
   sin[110]  =  16'b1101_1000_0000_0010;     //110pi/512
   cos[110]  =  16'b0011_0001_1111_0111;     //110pi/512
   sin[111]  =  16'b1101_0111_1011_0100;     //111pi/512
   cos[111]  =  16'b0011_0001_1011_1000;     //111pi/512
   sin[112]  =  16'b1101_0111_0110_0110;     //112pi/512
   cos[112]  =  16'b0011_0001_0111_1001;     //112pi/512
   sin[113]  =  16'b1101_0111_0001_1001;     //113pi/512
   cos[113]  =  16'b0011_0001_0011_1000;     //113pi/512
   sin[114]  =  16'b1101_0110_1100_1011;     //114pi/512
   cos[114]  =  16'b0011_0000_1111_1000;     //114pi/512
   sin[115]  =  16'b1101_0110_0111_1111;     //115pi/512
   cos[115]  =  16'b0011_0000_1011_0111;     //115pi/512
   sin[116]  =  16'b1101_0110_0011_0010;     //116pi/512
   cos[116]  =  16'b0011_0000_0111_0110;     //116pi/512
   sin[117]  =  16'b1101_0101_1110_0110;     //117pi/512
   cos[117]  =  16'b0011_0000_0011_0100;     //117pi/512
   sin[118]  =  16'b1101_0101_1001_1011;     //118pi/512
   cos[118]  =  16'b0010_1111_1111_0001;     //118pi/512
   sin[119]  =  16'b1101_0101_0101_0000;     //119pi/512
   cos[119]  =  16'b0010_1111_1010_1111;     //119pi/512
   sin[120]  =  16'b1101_0101_0000_0101;     //120pi/512
   cos[120]  =  16'b0010_1111_0110_1011;     //120pi/512
   sin[121]  =  16'b1101_0100_1011_1011;     //121pi/512
   cos[121]  =  16'b0010_1111_0010_1000;     //121pi/512
   sin[122]  =  16'b1101_0100_0111_0001;     //122pi/512
   cos[122]  =  16'b0010_1110_1110_0011;     //122pi/512
   sin[123]  =  16'b1101_0100_0010_1000;     //123pi/512
   cos[123]  =  16'b0010_1110_1001_1111;     //123pi/512
   sin[124]  =  16'b1101_0011_1101_1111;     //124pi/512
   cos[124]  =  16'b0010_1110_0101_1010;     //124pi/512
   sin[125]  =  16'b1101_0011_1001_0110;     //125pi/512
   cos[125]  =  16'b0010_1110_0001_0100;     //125pi/512
   sin[126]  =  16'b1101_0011_0100_1110;     //126pi/512
   cos[126]  =  16'b0010_1101_1100_1110;     //126pi/512
   sin[127]  =  16'b1101_0011_0000_0110;     //127pi/512
   cos[127]  =  16'b0010_1101_1000_1000;     //127pi/512
   sin[128]  =  16'b1101_0010_1011_1111;     //128pi/512
   cos[128]  =  16'b0010_1101_0100_0001;     //128pi/512
   sin[129]  =  16'b1101_0010_0111_1000;     //129pi/512
   cos[129]  =  16'b0010_1100_1111_1001;     //129pi/512
   sin[130]  =  16'b1101_0010_0011_0001;     //130pi/512
   cos[130]  =  16'b0010_1100_1011_0010;     //130pi/512
   sin[131]  =  16'b1101_0001_1110_1011;     //131pi/512
   cos[131]  =  16'b0010_1100_0110_1010;     //131pi/512
   sin[132]  =  16'b1101_0001_1010_0110;     //132pi/512
   cos[132]  =  16'b0010_1100_0010_0001;     //132pi/512
   sin[133]  =  16'b1101_0001_0110_0001;     //133pi/512
   cos[133]  =  16'b0010_1011_1101_1000;     //133pi/512
   sin[134]  =  16'b1101_0001_0001_1100;     //134pi/512
   cos[134]  =  16'b0010_1011_1000_1110;     //134pi/512
   sin[135]  =  16'b1101_0000_1101_1000;     //135pi/512
   cos[135]  =  16'b0010_1011_0100_0101;     //135pi/512
   sin[136]  =  16'b1101_0000_1001_0100;     //136pi/512
   cos[136]  =  16'b0010_1010_1111_1010;     //136pi/512
   sin[137]  =  16'b1101_0000_0101_0001;     //137pi/512
   cos[137]  =  16'b0010_1010_1011_0000;     //137pi/512
   sin[138]  =  16'b1101_0000_0000_1110;     //138pi/512
   cos[138]  =  16'b0010_1010_0110_0101;     //138pi/512
   sin[139]  =  16'b1100_1111_1100_1100;     //139pi/512
   cos[139]  =  16'b0010_1010_0001_1001;     //139pi/512
   sin[140]  =  16'b1100_1111_1000_1010;     //140pi/512
   cos[140]  =  16'b0010_1001_1100_1101;     //140pi/512
   sin[141]  =  16'b1100_1111_0100_1000;     //141pi/512
   cos[141]  =  16'b0010_1001_1000_0001;     //141pi/512
   sin[142]  =  16'b1100_1111_0000_0111;     //142pi/512
   cos[142]  =  16'b0010_1001_0011_0100;     //142pi/512
   sin[143]  =  16'b1100_1110_1100_0111;     //143pi/512
   cos[143]  =  16'b0010_1000_1110_0111;     //143pi/512
   sin[144]  =  16'b1100_1110_1000_0111;     //144pi/512
   cos[144]  =  16'b0010_1000_1001_1001;     //144pi/512
   sin[145]  =  16'b1100_1110_0100_0111;     //145pi/512
   cos[145]  =  16'b0010_1000_0100_1011;     //145pi/512
   sin[146]  =  16'b1100_1110_0000_1000;     //146pi/512
   cos[146]  =  16'b0010_0111_1111_1101;     //146pi/512
   sin[147]  =  16'b1100_1101_1100_1010;     //147pi/512
   cos[147]  =  16'b0010_0111_1010_1111;     //147pi/512
   sin[148]  =  16'b1100_1101_1000_1100;     //148pi/512
   cos[148]  =  16'b0010_0111_0101_1111;     //148pi/512
   sin[149]  =  16'b1100_1101_0100_1110;     //149pi/512
   cos[149]  =  16'b0010_0111_0001_0000;     //149pi/512
   sin[150]  =  16'b1100_1101_0001_0001;     //150pi/512
   cos[150]  =  16'b0010_0110_1100_0000;     //150pi/512
   sin[151]  =  16'b1100_1100_1101_0100;     //151pi/512
   cos[151]  =  16'b0010_0110_0111_0000;     //151pi/512
   sin[152]  =  16'b1100_1100_1001_1000;     //152pi/512
   cos[152]  =  16'b0010_0110_0001_1111;     //152pi/512
   sin[153]  =  16'b1100_1100_0101_1101;     //153pi/512
   cos[153]  =  16'b0010_0101_1100_1111;     //153pi/512
   sin[154]  =  16'b1100_1100_0010_0001;     //154pi/512
   cos[154]  =  16'b0010_0101_0111_1101;     //154pi/512
   sin[155]  =  16'b1100_1011_1110_0111;     //155pi/512
   cos[155]  =  16'b0010_0101_0010_1100;     //155pi/512
   sin[156]  =  16'b1100_1011_1010_1101;     //156pi/512
   cos[156]  =  16'b0010_0100_1101_1010;     //156pi/512
   sin[157]  =  16'b1100_1011_0111_0011;     //157pi/512
   cos[157]  =  16'b0010_0100_1000_0111;     //157pi/512
   sin[158]  =  16'b1100_1011_0011_1010;     //158pi/512
   cos[158]  =  16'b0010_0100_0011_0100;     //158pi/512
   sin[159]  =  16'b1100_1011_0000_0001;     //159pi/512
   cos[159]  =  16'b0010_0011_1110_0001;     //159pi/512
   sin[160]  =  16'b1100_1010_1100_1001;     //160pi/512
   cos[160]  =  16'b0010_0011_1000_1110;     //160pi/512
   sin[161]  =  16'b1100_1010_1001_0010;     //161pi/512
   cos[161]  =  16'b0010_0011_0011_1010;     //161pi/512
   sin[162]  =  16'b1100_1010_0101_1011;     //162pi/512
   cos[162]  =  16'b0010_0010_1110_0110;     //162pi/512
   sin[163]  =  16'b1100_1010_0010_0100;     //163pi/512
   cos[163]  =  16'b0010_0010_1001_0010;     //163pi/512
   sin[164]  =  16'b1100_1001_1110_1110;     //164pi/512
   cos[164]  =  16'b0010_0010_0011_1101;     //164pi/512
   sin[165]  =  16'b1100_1001_1011_1000;     //165pi/512
   cos[165]  =  16'b0010_0001_1110_1000;     //165pi/512
   sin[166]  =  16'b1100_1001_1000_0011;     //166pi/512
   cos[166]  =  16'b0010_0001_1001_0010;     //166pi/512
   sin[167]  =  16'b1100_1001_0100_1111;     //167pi/512
   cos[167]  =  16'b0010_0001_0011_1101;     //167pi/512
   sin[168]  =  16'b1100_1001_0001_1011;     //168pi/512
   cos[168]  =  16'b0010_0000_1110_0111;     //168pi/512
   sin[169]  =  16'b1100_1000_1110_1000;     //169pi/512
   cos[169]  =  16'b0010_0000_1001_0000;     //169pi/512
   sin[170]  =  16'b1100_1000_1011_0101;     //170pi/512
   cos[170]  =  16'b0010_0000_0011_1001;     //170pi/512
   sin[171]  =  16'b1100_1000_1000_0010;     //171pi/512
   cos[171]  =  16'b0001_1111_1110_0010;     //171pi/512
   sin[172]  =  16'b1100_1000_0101_0000;     //172pi/512
   cos[172]  =  16'b0001_1111_1000_1011;     //172pi/512
   sin[173]  =  16'b1100_1000_0001_1111;     //173pi/512
   cos[173]  =  16'b0001_1111_0011_0100;     //173pi/512
   sin[174]  =  16'b1100_0111_1110_1110;     //174pi/512
   cos[174]  =  16'b0001_1110_1101_1100;     //174pi/512
   sin[175]  =  16'b1100_0111_1011_1110;     //175pi/512
   cos[175]  =  16'b0001_1110_1000_0011;     //175pi/512
   sin[176]  =  16'b1100_0111_1000_1111;     //176pi/512
   cos[176]  =  16'b0001_1110_0010_1011;     //176pi/512
   sin[177]  =  16'b1100_0111_0101_1111;     //177pi/512
   cos[177]  =  16'b0001_1101_1101_0010;     //177pi/512
   sin[178]  =  16'b1100_0111_0011_0001;     //178pi/512
   cos[178]  =  16'b0001_1101_0111_1001;     //178pi/512
   sin[179]  =  16'b1100_0111_0000_0011;     //179pi/512
   cos[179]  =  16'b0001_1101_0010_0000;     //179pi/512
   sin[180]  =  16'b1100_0110_1101_0101;     //180pi/512
   cos[180]  =  16'b0001_1100_1100_0110;     //180pi/512
   sin[181]  =  16'b1100_0110_1010_1000;     //181pi/512
   cos[181]  =  16'b0001_1100_0110_1100;     //181pi/512
   sin[182]  =  16'b1100_0110_0111_1100;     //182pi/512
   cos[182]  =  16'b0001_1100_0001_0010;     //182pi/512
   sin[183]  =  16'b1100_0110_0101_0000;     //183pi/512
   cos[183]  =  16'b0001_1011_1011_0111;     //183pi/512
   sin[184]  =  16'b1100_0110_0010_0101;     //184pi/512
   cos[184]  =  16'b0001_1011_0101_1101;     //184pi/512
   sin[185]  =  16'b1100_0101_1111_1010;     //185pi/512
   cos[185]  =  16'b0001_1011_0000_0010;     //185pi/512
   sin[186]  =  16'b1100_0101_1101_0000;     //186pi/512
   cos[186]  =  16'b0001_1010_1010_0110;     //186pi/512
   sin[187]  =  16'b1100_0101_1010_0111;     //187pi/512
   cos[187]  =  16'b0001_1010_0100_1011;     //187pi/512
   sin[188]  =  16'b1100_0101_0111_1110;     //188pi/512
   cos[188]  =  16'b0001_1001_1110_1111;     //188pi/512
   sin[189]  =  16'b1100_0101_0101_0101;     //189pi/512
   cos[189]  =  16'b0001_1001_1001_0011;     //189pi/512
   sin[190]  =  16'b1100_0101_0010_1101;     //190pi/512
   cos[190]  =  16'b0001_1001_0011_0111;     //190pi/512
   sin[191]  =  16'b1100_0101_0000_0110;     //191pi/512
   cos[191]  =  16'b0001_1000_1101_1010;     //191pi/512
   sin[192]  =  16'b1100_0100_1101_1111;     //192pi/512
   cos[192]  =  16'b0001_1000_0111_1101;     //192pi/512
   sin[193]  =  16'b1100_0100_1011_1001;     //193pi/512
   cos[193]  =  16'b0001_1000_0010_0000;     //193pi/512
   sin[194]  =  16'b1100_0100_1001_0011;     //194pi/512
   cos[194]  =  16'b0001_0111_1100_0011;     //194pi/512
   sin[195]  =  16'b1100_0100_0110_1110;     //195pi/512
   cos[195]  =  16'b0001_0111_0110_0110;     //195pi/512
   sin[196]  =  16'b1100_0100_0100_1010;     //196pi/512
   cos[196]  =  16'b0001_0111_0000_1000;     //196pi/512
   sin[197]  =  16'b1100_0100_0010_0110;     //197pi/512
   cos[197]  =  16'b0001_0110_1010_1010;     //197pi/512
   sin[198]  =  16'b1100_0100_0000_0011;     //198pi/512
   cos[198]  =  16'b0001_0110_0100_1100;     //198pi/512
   sin[199]  =  16'b1100_0011_1110_0000;     //199pi/512
   cos[199]  =  16'b0001_0101_1110_1110;     //199pi/512
   sin[200]  =  16'b1100_0011_1011_1110;     //200pi/512
   cos[200]  =  16'b0001_0101_1000_1111;     //200pi/512
   sin[201]  =  16'b1100_0011_1001_1100;     //201pi/512
   cos[201]  =  16'b0001_0101_0011_0000;     //201pi/512
   sin[202]  =  16'b1100_0011_0111_1011;     //202pi/512
   cos[202]  =  16'b0001_0100_1101_0001;     //202pi/512
   sin[203]  =  16'b1100_0011_0101_1011;     //203pi/512
   cos[203]  =  16'b0001_0100_0111_0010;     //203pi/512
   sin[204]  =  16'b1100_0011_0011_1011;     //204pi/512
   cos[204]  =  16'b0001_0100_0001_0011;     //204pi/512
   sin[205]  =  16'b1100_0011_0001_1100;     //205pi/512
   cos[205]  =  16'b0001_0011_1011_0011;     //205pi/512
   sin[206]  =  16'b1100_0010_1111_1101;     //206pi/512
   cos[206]  =  16'b0001_0011_0101_0100;     //206pi/512
   sin[207]  =  16'b1100_0010_1101_1111;     //207pi/512
   cos[207]  =  16'b0001_0010_1111_0100;     //207pi/512
   sin[208]  =  16'b1100_0010_1100_0001;     //208pi/512
   cos[208]  =  16'b0001_0010_1001_0100;     //208pi/512
   sin[209]  =  16'b1100_0010_1010_0101;     //209pi/512
   cos[209]  =  16'b0001_0010_0011_0011;     //209pi/512
   sin[210]  =  16'b1100_0010_1000_1000;     //210pi/512
   cos[210]  =  16'b0001_0001_1101_0011;     //210pi/512
   sin[211]  =  16'b1100_0010_0110_1101;     //211pi/512
   cos[211]  =  16'b0001_0001_0111_0010;     //211pi/512
   sin[212]  =  16'b1100_0010_0101_0001;     //212pi/512
   cos[212]  =  16'b0001_0001_0001_0001;     //212pi/512
   sin[213]  =  16'b1100_0010_0011_0111;     //213pi/512
   cos[213]  =  16'b0001_0000_1011_0000;     //213pi/512
   sin[214]  =  16'b1100_0010_0001_1101;     //214pi/512
   cos[214]  =  16'b0001_0000_0100_1111;     //214pi/512
   sin[215]  =  16'b1100_0010_0000_0100;     //215pi/512
   cos[215]  =  16'b0000_1111_1110_1110;     //215pi/512
   sin[216]  =  16'b1100_0001_1110_1011;     //216pi/512
   cos[216]  =  16'b0000_1111_1000_1100;     //216pi/512
   sin[217]  =  16'b1100_0001_1101_0011;     //217pi/512
   cos[217]  =  16'b0000_1111_0010_1011;     //217pi/512
   sin[218]  =  16'b1100_0001_1011_1011;     //218pi/512
   cos[218]  =  16'b0000_1110_1100_1001;     //218pi/512
   sin[219]  =  16'b1100_0001_1010_0100;     //219pi/512
   cos[219]  =  16'b0000_1110_0110_0111;     //219pi/512
   sin[220]  =  16'b1100_0001_1000_1110;     //220pi/512
   cos[220]  =  16'b0000_1110_0000_0101;     //220pi/512
   sin[221]  =  16'b1100_0001_0111_1000;     //221pi/512
   cos[221]  =  16'b0000_1101_1010_0011;     //221pi/512
   sin[222]  =  16'b1100_0001_0110_0011;     //222pi/512
   cos[222]  =  16'b0000_1101_0100_0001;     //222pi/512
   sin[223]  =  16'b1100_0001_0100_1111;     //223pi/512
   cos[223]  =  16'b0000_1100_1101_1110;     //223pi/512
   sin[224]  =  16'b1100_0001_0011_1011;     //224pi/512
   cos[224]  =  16'b0000_1100_0111_1100;     //224pi/512
   sin[225]  =  16'b1100_0001_0010_1000;     //225pi/512
   cos[225]  =  16'b0000_1100_0001_1001;     //225pi/512
   sin[226]  =  16'b1100_0001_0001_0101;     //226pi/512
   cos[226]  =  16'b0000_1011_1011_0110;     //226pi/512
   sin[227]  =  16'b1100_0001_0000_0011;     //227pi/512
   cos[227]  =  16'b0000_1011_0101_0100;     //227pi/512
   sin[228]  =  16'b1100_0000_1111_0001;     //228pi/512
   cos[228]  =  16'b0000_1010_1111_0001;     //228pi/512
   sin[229]  =  16'b1100_0000_1110_0000;     //229pi/512
   cos[229]  =  16'b0000_1010_1000_1101;     //229pi/512
   sin[230]  =  16'b1100_0000_1101_0000;     //230pi/512
   cos[230]  =  16'b0000_1010_0010_1010;     //230pi/512
   sin[231]  =  16'b1100_0000_1100_0000;     //231pi/512
   cos[231]  =  16'b0000_1001_1100_0111;     //231pi/512
   sin[232]  =  16'b1100_0000_1011_0001;     //232pi/512
   cos[232]  =  16'b0000_1001_0110_0100;     //232pi/512
   sin[233]  =  16'b1100_0000_1010_0011;     //233pi/512
   cos[233]  =  16'b0000_1001_0000_0000;     //233pi/512
   sin[234]  =  16'b1100_0000_1001_0101;     //234pi/512
   cos[234]  =  16'b0000_1000_1001_1100;     //234pi/512
   sin[235]  =  16'b1100_0000_1000_1000;     //235pi/512
   cos[235]  =  16'b0000_1000_0011_1001;     //235pi/512
   sin[236]  =  16'b1100_0000_0111_1011;     //236pi/512
   cos[236]  =  16'b0000_0111_1101_0101;     //236pi/512
   sin[237]  =  16'b1100_0000_0110_1111;     //237pi/512
   cos[237]  =  16'b0000_0111_0111_0001;     //237pi/512
   sin[238]  =  16'b1100_0000_0110_0100;     //238pi/512
   cos[238]  =  16'b0000_0111_0000_1101;     //238pi/512
   sin[239]  =  16'b1100_0000_0101_1001;     //239pi/512
   cos[239]  =  16'b0000_0110_1010_1001;     //239pi/512
   sin[240]  =  16'b1100_0000_0100_1111;     //240pi/512
   cos[240]  =  16'b0000_0110_0100_0101;     //240pi/512
   sin[241]  =  16'b1100_0000_0100_0101;     //241pi/512
   cos[241]  =  16'b0000_0101_1110_0001;     //241pi/512
   sin[242]  =  16'b1100_0000_0011_1100;     //242pi/512
   cos[242]  =  16'b0000_0101_0111_1101;     //242pi/512
   sin[243]  =  16'b1100_0000_0011_0100;     //243pi/512
   cos[243]  =  16'b0000_0101_0001_1001;     //243pi/512
   sin[244]  =  16'b1100_0000_0010_1100;     //244pi/512
   cos[244]  =  16'b0000_0100_1011_0101;     //244pi/512
   sin[245]  =  16'b1100_0000_0010_0101;     //245pi/512
   cos[245]  =  16'b0000_0100_0101_0001;     //245pi/512
   sin[246]  =  16'b1100_0000_0001_1111;     //246pi/512
   cos[246]  =  16'b0000_0011_1110_1100;     //246pi/512
   sin[247]  =  16'b1100_0000_0001_1001;     //247pi/512
   cos[247]  =  16'b0000_0011_1000_1000;     //247pi/512
   sin[248]  =  16'b1100_0000_0001_0100;     //248pi/512
   cos[248]  =  16'b0000_0011_0010_0011;     //248pi/512
   sin[249]  =  16'b1100_0000_0000_1111;     //249pi/512
   cos[249]  =  16'b0000_0010_1011_1111;     //249pi/512
   sin[250]  =  16'b1100_0000_0000_1011;     //250pi/512
   cos[250]  =  16'b0000_0010_0101_1011;     //250pi/512
   sin[251]  =  16'b1100_0000_0000_1000;     //251pi/512
   cos[251]  =  16'b0000_0001_1111_0110;     //251pi/512
   sin[252]  =  16'b1100_0000_0000_0101;     //252pi/512
   cos[252]  =  16'b0000_0001_1001_0010;     //252pi/512
   sin[253]  =  16'b1100_0000_0000_0011;     //253pi/512
   cos[253]  =  16'b0000_0001_0010_1101;     //253pi/512
   sin[254]  =  16'b1100_0000_0000_0001;     //254pi/512
   cos[254]  =  16'b0000_0000_1100_1001;     //254pi/512
   sin[255]  =  16'b1100_0000_0000_0000;     //255pi/512
   cos[255]  =  16'b0000_0000_0110_0100;     //255pi/512
   sin[256]  =  16'b1100_0000_0000_0000;     //256pi/512
   cos[256]  =  16'b0000_0000_0000_0000;     //256pi/512
   sin[257]  =  16'b1100_0000_0000_0000;     //257pi/512
   cos[257]  =  16'b1111_1111_1001_1011;     //257pi/512
   sin[258]  =  16'b1100_0000_0000_0001;     //258pi/512
   cos[258]  =  16'b1111_1111_0011_0111;     //258pi/512
   sin[259]  =  16'b1100_0000_0000_0011;     //259pi/512
   cos[259]  =  16'b1111_1110_1101_0010;     //259pi/512
   sin[260]  =  16'b1100_0000_0000_0101;     //260pi/512
   cos[260]  =  16'b1111_1110_0110_1110;     //260pi/512
   sin[261]  =  16'b1100_0000_0000_1000;     //261pi/512
   cos[261]  =  16'b1111_1110_0000_1001;     //261pi/512
   sin[262]  =  16'b1100_0000_0000_1011;     //262pi/512
   cos[262]  =  16'b1111_1101_1010_0101;     //262pi/512
   sin[263]  =  16'b1100_0000_0000_1111;     //263pi/512
   cos[263]  =  16'b1111_1101_0100_0000;     //263pi/512
   sin[264]  =  16'b1100_0000_0001_0100;     //264pi/512
   cos[264]  =  16'b1111_1100_1101_1100;     //264pi/512
   sin[265]  =  16'b1100_0000_0001_1001;     //265pi/512
   cos[265]  =  16'b1111_1100_0111_1000;     //265pi/512
   sin[266]  =  16'b1100_0000_0001_1111;     //266pi/512
   cos[266]  =  16'b1111_1100_0001_0011;     //266pi/512
   sin[267]  =  16'b1100_0000_0010_0101;     //267pi/512
   cos[267]  =  16'b1111_1011_1010_1111;     //267pi/512
   sin[268]  =  16'b1100_0000_0010_1100;     //268pi/512
   cos[268]  =  16'b1111_1011_0100_1011;     //268pi/512
   sin[269]  =  16'b1100_0000_0011_0100;     //269pi/512
   cos[269]  =  16'b1111_1010_1110_0110;     //269pi/512
   sin[270]  =  16'b1100_0000_0011_1100;     //270pi/512
   cos[270]  =  16'b1111_1010_1000_0010;     //270pi/512
   sin[271]  =  16'b1100_0000_0100_0101;     //271pi/512
   cos[271]  =  16'b1111_1010_0001_1110;     //271pi/512
   sin[272]  =  16'b1100_0000_0100_1111;     //272pi/512
   cos[272]  =  16'b1111_1001_1011_1010;     //272pi/512
   sin[273]  =  16'b1100_0000_0101_1001;     //273pi/512
   cos[273]  =  16'b1111_1001_0101_0110;     //273pi/512
   sin[274]  =  16'b1100_0000_0110_0100;     //274pi/512
   cos[274]  =  16'b1111_1000_1111_0010;     //274pi/512
   sin[275]  =  16'b1100_0000_0110_1111;     //275pi/512
   cos[275]  =  16'b1111_1000_1000_1110;     //275pi/512
   sin[276]  =  16'b1100_0000_0111_1011;     //276pi/512
   cos[276]  =  16'b1111_1000_0010_1010;     //276pi/512
   sin[277]  =  16'b1100_0000_1000_1000;     //277pi/512
   cos[277]  =  16'b1111_0111_1100_0111;     //277pi/512
   sin[278]  =  16'b1100_0000_1001_0101;     //278pi/512
   cos[278]  =  16'b1111_0111_0110_0011;     //278pi/512
   sin[279]  =  16'b1100_0000_1010_0011;     //279pi/512
   cos[279]  =  16'b1111_0110_1111_1111;     //279pi/512
   sin[280]  =  16'b1100_0000_1011_0001;     //280pi/512
   cos[280]  =  16'b1111_0110_1001_1100;     //280pi/512
   sin[281]  =  16'b1100_0000_1100_0000;     //281pi/512
   cos[281]  =  16'b1111_0110_0011_1001;     //281pi/512
   sin[282]  =  16'b1100_0000_1101_0000;     //282pi/512
   cos[282]  =  16'b1111_0101_1101_0101;     //282pi/512
   sin[283]  =  16'b1100_0000_1110_0000;     //283pi/512
   cos[283]  =  16'b1111_0101_0111_0010;     //283pi/512
   sin[284]  =  16'b1100_0000_1111_0001;     //284pi/512
   cos[284]  =  16'b1111_0101_0000_1111;     //284pi/512
   sin[285]  =  16'b1100_0001_0000_0011;     //285pi/512
   cos[285]  =  16'b1111_0100_1010_1100;     //285pi/512
   sin[286]  =  16'b1100_0001_0001_0101;     //286pi/512
   cos[286]  =  16'b1111_0100_0100_1001;     //286pi/512
   sin[287]  =  16'b1100_0001_0010_1000;     //287pi/512
   cos[287]  =  16'b1111_0011_1110_0110;     //287pi/512
   sin[288]  =  16'b1100_0001_0011_1011;     //288pi/512
   cos[288]  =  16'b1111_0011_1000_0100;     //288pi/512
   sin[289]  =  16'b1100_0001_0100_1111;     //289pi/512
   cos[289]  =  16'b1111_0011_0010_0001;     //289pi/512
   sin[290]  =  16'b1100_0001_0110_0011;     //290pi/512
   cos[290]  =  16'b1111_0010_1011_1111;     //290pi/512
   sin[291]  =  16'b1100_0001_0111_1000;     //291pi/512
   cos[291]  =  16'b1111_0010_0101_1100;     //291pi/512
   sin[292]  =  16'b1100_0001_1000_1110;     //292pi/512
   cos[292]  =  16'b1111_0001_1111_1010;     //292pi/512
   sin[293]  =  16'b1100_0001_1010_0100;     //293pi/512
   cos[293]  =  16'b1111_0001_1001_1000;     //293pi/512
   sin[294]  =  16'b1100_0001_1011_1011;     //294pi/512
   cos[294]  =  16'b1111_0001_0011_0110;     //294pi/512
   sin[295]  =  16'b1100_0001_1101_0011;     //295pi/512
   cos[295]  =  16'b1111_0000_1101_0101;     //295pi/512
   sin[296]  =  16'b1100_0001_1110_1011;     //296pi/512
   cos[296]  =  16'b1111_0000_0111_0011;     //296pi/512
   sin[297]  =  16'b1100_0010_0000_0100;     //297pi/512
   cos[297]  =  16'b1111_0000_0001_0010;     //297pi/512
   sin[298]  =  16'b1100_0010_0001_1101;     //298pi/512
   cos[298]  =  16'b1110_1111_1011_0000;     //298pi/512
   sin[299]  =  16'b1100_0010_0011_0111;     //299pi/512
   cos[299]  =  16'b1110_1111_0100_1111;     //299pi/512
   sin[300]  =  16'b1100_0010_0101_0001;     //300pi/512
   cos[300]  =  16'b1110_1110_1110_1110;     //300pi/512
   sin[301]  =  16'b1100_0010_0110_1101;     //301pi/512
   cos[301]  =  16'b1110_1110_1000_1101;     //301pi/512
   sin[302]  =  16'b1100_0010_1000_1000;     //302pi/512
   cos[302]  =  16'b1110_1110_0010_1101;     //302pi/512
   sin[303]  =  16'b1100_0010_1010_0101;     //303pi/512
   cos[303]  =  16'b1110_1101_1100_1100;     //303pi/512
   sin[304]  =  16'b1100_0010_1100_0001;     //304pi/512
   cos[304]  =  16'b1110_1101_0110_1100;     //304pi/512
   sin[305]  =  16'b1100_0010_1101_1111;     //305pi/512
   cos[305]  =  16'b1110_1101_0000_1100;     //305pi/512
   sin[306]  =  16'b1100_0010_1111_1101;     //306pi/512
   cos[306]  =  16'b1110_1100_1010_1100;     //306pi/512
   sin[307]  =  16'b1100_0011_0001_1100;     //307pi/512
   cos[307]  =  16'b1110_1100_0100_1100;     //307pi/512
   sin[308]  =  16'b1100_0011_0011_1011;     //308pi/512
   cos[308]  =  16'b1110_1011_1110_1101;     //308pi/512
   sin[309]  =  16'b1100_0011_0101_1011;     //309pi/512
   cos[309]  =  16'b1110_1011_1000_1101;     //309pi/512
   sin[310]  =  16'b1100_0011_0111_1011;     //310pi/512
   cos[310]  =  16'b1110_1011_0010_1110;     //310pi/512
   sin[311]  =  16'b1100_0011_1001_1100;     //311pi/512
   cos[311]  =  16'b1110_1010_1100_1111;     //311pi/512
   sin[312]  =  16'b1100_0011_1011_1110;     //312pi/512
   cos[312]  =  16'b1110_1010_0111_0000;     //312pi/512
   sin[313]  =  16'b1100_0011_1110_0000;     //313pi/512
   cos[313]  =  16'b1110_1010_0001_0010;     //313pi/512
   sin[314]  =  16'b1100_0100_0000_0011;     //314pi/512
   cos[314]  =  16'b1110_1001_1011_0100;     //314pi/512
   sin[315]  =  16'b1100_0100_0010_0110;     //315pi/512
   cos[315]  =  16'b1110_1001_0101_0101;     //315pi/512
   sin[316]  =  16'b1100_0100_0100_1010;     //316pi/512
   cos[316]  =  16'b1110_1000_1111_0111;     //316pi/512
   sin[317]  =  16'b1100_0100_0110_1110;     //317pi/512
   cos[317]  =  16'b1110_1000_1001_1010;     //317pi/512
   sin[318]  =  16'b1100_0100_1001_0011;     //318pi/512
   cos[318]  =  16'b1110_1000_0011_1100;     //318pi/512
   sin[319]  =  16'b1100_0100_1011_1001;     //319pi/512
   cos[319]  =  16'b1110_0111_1101_1111;     //319pi/512
   sin[320]  =  16'b1100_0100_1101_1111;     //320pi/512
   cos[320]  =  16'b1110_0111_1000_0010;     //320pi/512
   sin[321]  =  16'b1100_0101_0000_0110;     //321pi/512
   cos[321]  =  16'b1110_0111_0010_0101;     //321pi/512
   sin[322]  =  16'b1100_0101_0010_1101;     //322pi/512
   cos[322]  =  16'b1110_0110_1100_1001;     //322pi/512
   sin[323]  =  16'b1100_0101_0101_0101;     //323pi/512
   cos[323]  =  16'b1110_0110_0110_1101;     //323pi/512
   sin[324]  =  16'b1100_0101_0111_1110;     //324pi/512
   cos[324]  =  16'b1110_0110_0001_0001;     //324pi/512
   sin[325]  =  16'b1100_0101_1010_0111;     //325pi/512
   cos[325]  =  16'b1110_0101_1011_0101;     //325pi/512
   sin[326]  =  16'b1100_0101_1101_0000;     //326pi/512
   cos[326]  =  16'b1110_0101_0101_1001;     //326pi/512
   sin[327]  =  16'b1100_0101_1111_1010;     //327pi/512
   cos[327]  =  16'b1110_0100_1111_1110;     //327pi/512
   sin[328]  =  16'b1100_0110_0010_0101;     //328pi/512
   cos[328]  =  16'b1110_0100_1010_0011;     //328pi/512
   sin[329]  =  16'b1100_0110_0101_0000;     //329pi/512
   cos[329]  =  16'b1110_0100_0100_1000;     //329pi/512
   sin[330]  =  16'b1100_0110_0111_1100;     //330pi/512
   cos[330]  =  16'b1110_0011_1110_1110;     //330pi/512
   sin[331]  =  16'b1100_0110_1010_1000;     //331pi/512
   cos[331]  =  16'b1110_0011_1001_0100;     //331pi/512
   sin[332]  =  16'b1100_0110_1101_0101;     //332pi/512
   cos[332]  =  16'b1110_0011_0011_1010;     //332pi/512
   sin[333]  =  16'b1100_0111_0000_0011;     //333pi/512
   cos[333]  =  16'b1110_0010_1110_0000;     //333pi/512
   sin[334]  =  16'b1100_0111_0011_0001;     //334pi/512
   cos[334]  =  16'b1110_0010_1000_0111;     //334pi/512
   sin[335]  =  16'b1100_0111_0101_1111;     //335pi/512
   cos[335]  =  16'b1110_0010_0010_1101;     //335pi/512
   sin[336]  =  16'b1100_0111_1000_1111;     //336pi/512
   cos[336]  =  16'b1110_0001_1101_0101;     //336pi/512
   sin[337]  =  16'b1100_0111_1011_1110;     //337pi/512
   cos[337]  =  16'b1110_0001_0111_1100;     //337pi/512
   sin[338]  =  16'b1100_0111_1110_1110;     //338pi/512
   cos[338]  =  16'b1110_0001_0010_0100;     //338pi/512
   sin[339]  =  16'b1100_1000_0001_1111;     //339pi/512
   cos[339]  =  16'b1110_0000_1100_1100;     //339pi/512
   sin[340]  =  16'b1100_1000_0101_0000;     //340pi/512
   cos[340]  =  16'b1110_0000_0111_0100;     //340pi/512
   sin[341]  =  16'b1100_1000_1000_0010;     //341pi/512
   cos[341]  =  16'b1110_0000_0001_1101;     //341pi/512
   sin[342]  =  16'b1100_1000_1011_0101;     //342pi/512
   cos[342]  =  16'b1101_1111_1100_0110;     //342pi/512
   sin[343]  =  16'b1100_1000_1110_1000;     //343pi/512
   cos[343]  =  16'b1101_1111_0110_1111;     //343pi/512
   sin[344]  =  16'b1100_1001_0001_1011;     //344pi/512
   cos[344]  =  16'b1101_1111_0001_1001;     //344pi/512
   sin[345]  =  16'b1100_1001_0100_1111;     //345pi/512
   cos[345]  =  16'b1101_1110_1100_0011;     //345pi/512
   sin[346]  =  16'b1100_1001_1000_0011;     //346pi/512
   cos[346]  =  16'b1101_1110_0110_1101;     //346pi/512
   sin[347]  =  16'b1100_1001_1011_1000;     //347pi/512
   cos[347]  =  16'b1101_1110_0001_1000;     //347pi/512
   sin[348]  =  16'b1100_1001_1110_1110;     //348pi/512
   cos[348]  =  16'b1101_1101_1100_0011;     //348pi/512
   sin[349]  =  16'b1100_1010_0010_0100;     //349pi/512
   cos[349]  =  16'b1101_1101_0110_1110;     //349pi/512
   sin[350]  =  16'b1100_1010_0101_1011;     //350pi/512
   cos[350]  =  16'b1101_1101_0001_1001;     //350pi/512
   sin[351]  =  16'b1100_1010_1001_0010;     //351pi/512
   cos[351]  =  16'b1101_1100_1100_0101;     //351pi/512
   sin[352]  =  16'b1100_1010_1100_1001;     //352pi/512
   cos[352]  =  16'b1101_1100_0111_0010;     //352pi/512
   sin[353]  =  16'b1100_1011_0000_0001;     //353pi/512
   cos[353]  =  16'b1101_1100_0001_1110;     //353pi/512
   sin[354]  =  16'b1100_1011_0011_1010;     //354pi/512
   cos[354]  =  16'b1101_1011_1100_1011;     //354pi/512
   sin[355]  =  16'b1100_1011_0111_0011;     //355pi/512
   cos[355]  =  16'b1101_1011_0111_1000;     //355pi/512
   sin[356]  =  16'b1100_1011_1010_1101;     //356pi/512
   cos[356]  =  16'b1101_1011_0010_0110;     //356pi/512
   sin[357]  =  16'b1100_1011_1110_0111;     //357pi/512
   cos[357]  =  16'b1101_1010_1101_0100;     //357pi/512
   sin[358]  =  16'b1100_1100_0010_0001;     //358pi/512
   cos[358]  =  16'b1101_1010_1000_0010;     //358pi/512
   sin[359]  =  16'b1100_1100_0101_1101;     //359pi/512
   cos[359]  =  16'b1101_1010_0011_0001;     //359pi/512
   sin[360]  =  16'b1100_1100_1001_1000;     //360pi/512
   cos[360]  =  16'b1101_1001_1110_0000;     //360pi/512
   sin[361]  =  16'b1100_1100_1101_0100;     //361pi/512
   cos[361]  =  16'b1101_1001_1000_1111;     //361pi/512
   sin[362]  =  16'b1100_1101_0001_0001;     //362pi/512
   cos[362]  =  16'b1101_1001_0011_1111;     //362pi/512
   sin[363]  =  16'b1100_1101_0100_1110;     //363pi/512
   cos[363]  =  16'b1101_1000_1110_1111;     //363pi/512
   sin[364]  =  16'b1100_1101_1000_1100;     //364pi/512
   cos[364]  =  16'b1101_1000_1010_0000;     //364pi/512
   sin[365]  =  16'b1100_1101_1100_1010;     //365pi/512
   cos[365]  =  16'b1101_1000_0101_0001;     //365pi/512
   sin[366]  =  16'b1100_1110_0000_1000;     //366pi/512
   cos[366]  =  16'b1101_1000_0000_0010;     //366pi/512
   sin[367]  =  16'b1100_1110_0100_0111;     //367pi/512
   cos[367]  =  16'b1101_0111_1011_0100;     //367pi/512
   sin[368]  =  16'b1100_1110_1000_0111;     //368pi/512
   cos[368]  =  16'b1101_0111_0110_0110;     //368pi/512
   sin[369]  =  16'b1100_1110_1100_0111;     //369pi/512
   cos[369]  =  16'b1101_0111_0001_1001;     //369pi/512
   sin[370]  =  16'b1100_1111_0000_0111;     //370pi/512
   cos[370]  =  16'b1101_0110_1100_1011;     //370pi/512
   sin[371]  =  16'b1100_1111_0100_1000;     //371pi/512
   cos[371]  =  16'b1101_0110_0111_1111;     //371pi/512
   sin[372]  =  16'b1100_1111_1000_1010;     //372pi/512
   cos[372]  =  16'b1101_0110_0011_0010;     //372pi/512
   sin[373]  =  16'b1100_1111_1100_1100;     //373pi/512
   cos[373]  =  16'b1101_0101_1110_0110;     //373pi/512
   sin[374]  =  16'b1101_0000_0000_1110;     //374pi/512
   cos[374]  =  16'b1101_0101_1001_1011;     //374pi/512
   sin[375]  =  16'b1101_0000_0101_0001;     //375pi/512
   cos[375]  =  16'b1101_0101_0101_0000;     //375pi/512
   sin[376]  =  16'b1101_0000_1001_0100;     //376pi/512
   cos[376]  =  16'b1101_0101_0000_0101;     //376pi/512
   sin[377]  =  16'b1101_0000_1101_1000;     //377pi/512
   cos[377]  =  16'b1101_0100_1011_1011;     //377pi/512
   sin[378]  =  16'b1101_0001_0001_1100;     //378pi/512
   cos[378]  =  16'b1101_0100_0111_0001;     //378pi/512
   sin[379]  =  16'b1101_0001_0110_0001;     //379pi/512
   cos[379]  =  16'b1101_0100_0010_1000;     //379pi/512
   sin[380]  =  16'b1101_0001_1010_0110;     //380pi/512
   cos[380]  =  16'b1101_0011_1101_1111;     //380pi/512
   sin[381]  =  16'b1101_0001_1110_1011;     //381pi/512
   cos[381]  =  16'b1101_0011_1001_0110;     //381pi/512
   sin[382]  =  16'b1101_0010_0011_0001;     //382pi/512
   cos[382]  =  16'b1101_0011_0100_1110;     //382pi/512
   sin[383]  =  16'b1101_0010_0111_1000;     //383pi/512
   cos[383]  =  16'b1101_0011_0000_0110;     //383pi/512
   sin[384]  =  16'b1101_0010_1011_1111;     //384pi/512
   cos[384]  =  16'b1101_0010_1011_1111;     //384pi/512
   sin[385]  =  16'b1101_0011_0000_0110;     //385pi/512
   cos[385]  =  16'b1101_0010_0111_1000;     //385pi/512
   sin[386]  =  16'b1101_0011_0100_1110;     //386pi/512
   cos[386]  =  16'b1101_0010_0011_0001;     //386pi/512
   sin[387]  =  16'b1101_0011_1001_0110;     //387pi/512
   cos[387]  =  16'b1101_0001_1110_1011;     //387pi/512
   sin[388]  =  16'b1101_0011_1101_1111;     //388pi/512
   cos[388]  =  16'b1101_0001_1010_0110;     //388pi/512
   sin[389]  =  16'b1101_0100_0010_1000;     //389pi/512
   cos[389]  =  16'b1101_0001_0110_0001;     //389pi/512
   sin[390]  =  16'b1101_0100_0111_0001;     //390pi/512
   cos[390]  =  16'b1101_0001_0001_1100;     //390pi/512
   sin[391]  =  16'b1101_0100_1011_1011;     //391pi/512
   cos[391]  =  16'b1101_0000_1101_1000;     //391pi/512
   sin[392]  =  16'b1101_0101_0000_0101;     //392pi/512
   cos[392]  =  16'b1101_0000_1001_0100;     //392pi/512
   sin[393]  =  16'b1101_0101_0101_0000;     //393pi/512
   cos[393]  =  16'b1101_0000_0101_0001;     //393pi/512
   sin[394]  =  16'b1101_0101_1001_1011;     //394pi/512
   cos[394]  =  16'b1101_0000_0000_1110;     //394pi/512
   sin[395]  =  16'b1101_0101_1110_0110;     //395pi/512
   cos[395]  =  16'b1100_1111_1100_1100;     //395pi/512
   sin[396]  =  16'b1101_0110_0011_0010;     //396pi/512
   cos[396]  =  16'b1100_1111_1000_1010;     //396pi/512
   sin[397]  =  16'b1101_0110_0111_1111;     //397pi/512
   cos[397]  =  16'b1100_1111_0100_1000;     //397pi/512
   sin[398]  =  16'b1101_0110_1100_1011;     //398pi/512
   cos[398]  =  16'b1100_1111_0000_0111;     //398pi/512
   sin[399]  =  16'b1101_0111_0001_1001;     //399pi/512
   cos[399]  =  16'b1100_1110_1100_0111;     //399pi/512
   sin[400]  =  16'b1101_0111_0110_0110;     //400pi/512
   cos[400]  =  16'b1100_1110_1000_0111;     //400pi/512
   sin[401]  =  16'b1101_0111_1011_0100;     //401pi/512
   cos[401]  =  16'b1100_1110_0100_0111;     //401pi/512
   sin[402]  =  16'b1101_1000_0000_0010;     //402pi/512
   cos[402]  =  16'b1100_1110_0000_1000;     //402pi/512
   sin[403]  =  16'b1101_1000_0101_0001;     //403pi/512
   cos[403]  =  16'b1100_1101_1100_1010;     //403pi/512
   sin[404]  =  16'b1101_1000_1010_0000;     //404pi/512
   cos[404]  =  16'b1100_1101_1000_1100;     //404pi/512
   sin[405]  =  16'b1101_1000_1110_1111;     //405pi/512
   cos[405]  =  16'b1100_1101_0100_1110;     //405pi/512
   sin[406]  =  16'b1101_1001_0011_1111;     //406pi/512
   cos[406]  =  16'b1100_1101_0001_0001;     //406pi/512
   sin[407]  =  16'b1101_1001_1000_1111;     //407pi/512
   cos[407]  =  16'b1100_1100_1101_0100;     //407pi/512
   sin[408]  =  16'b1101_1001_1110_0000;     //408pi/512
   cos[408]  =  16'b1100_1100_1001_1000;     //408pi/512
   sin[409]  =  16'b1101_1010_0011_0001;     //409pi/512
   cos[409]  =  16'b1100_1100_0101_1101;     //409pi/512
   sin[410]  =  16'b1101_1010_1000_0010;     //410pi/512
   cos[410]  =  16'b1100_1100_0010_0001;     //410pi/512
   sin[411]  =  16'b1101_1010_1101_0100;     //411pi/512
   cos[411]  =  16'b1100_1011_1110_0111;     //411pi/512
   sin[412]  =  16'b1101_1011_0010_0110;     //412pi/512
   cos[412]  =  16'b1100_1011_1010_1101;     //412pi/512
   sin[413]  =  16'b1101_1011_0111_1000;     //413pi/512
   cos[413]  =  16'b1100_1011_0111_0011;     //413pi/512
   sin[414]  =  16'b1101_1011_1100_1011;     //414pi/512
   cos[414]  =  16'b1100_1011_0011_1010;     //414pi/512
   sin[415]  =  16'b1101_1100_0001_1110;     //415pi/512
   cos[415]  =  16'b1100_1011_0000_0001;     //415pi/512
   sin[416]  =  16'b1101_1100_0111_0010;     //416pi/512
   cos[416]  =  16'b1100_1010_1100_1001;     //416pi/512
   sin[417]  =  16'b1101_1100_1100_0101;     //417pi/512
   cos[417]  =  16'b1100_1010_1001_0010;     //417pi/512
   sin[418]  =  16'b1101_1101_0001_1001;     //418pi/512
   cos[418]  =  16'b1100_1010_0101_1011;     //418pi/512
   sin[419]  =  16'b1101_1101_0110_1110;     //419pi/512
   cos[419]  =  16'b1100_1010_0010_0100;     //419pi/512
   sin[420]  =  16'b1101_1101_1100_0011;     //420pi/512
   cos[420]  =  16'b1100_1001_1110_1110;     //420pi/512
   sin[421]  =  16'b1101_1110_0001_1000;     //421pi/512
   cos[421]  =  16'b1100_1001_1011_1000;     //421pi/512
   sin[422]  =  16'b1101_1110_0110_1101;     //422pi/512
   cos[422]  =  16'b1100_1001_1000_0011;     //422pi/512
   sin[423]  =  16'b1101_1110_1100_0011;     //423pi/512
   cos[423]  =  16'b1100_1001_0100_1111;     //423pi/512
   sin[424]  =  16'b1101_1111_0001_1001;     //424pi/512
   cos[424]  =  16'b1100_1001_0001_1011;     //424pi/512
   sin[425]  =  16'b1101_1111_0110_1111;     //425pi/512
   cos[425]  =  16'b1100_1000_1110_1000;     //425pi/512
   sin[426]  =  16'b1101_1111_1100_0110;     //426pi/512
   cos[426]  =  16'b1100_1000_1011_0101;     //426pi/512
   sin[427]  =  16'b1110_0000_0001_1101;     //427pi/512
   cos[427]  =  16'b1100_1000_1000_0010;     //427pi/512
   sin[428]  =  16'b1110_0000_0111_0100;     //428pi/512
   cos[428]  =  16'b1100_1000_0101_0000;     //428pi/512
   sin[429]  =  16'b1110_0000_1100_1100;     //429pi/512
   cos[429]  =  16'b1100_1000_0001_1111;     //429pi/512
   sin[430]  =  16'b1110_0001_0010_0100;     //430pi/512
   cos[430]  =  16'b1100_0111_1110_1110;     //430pi/512
   sin[431]  =  16'b1110_0001_0111_1100;     //431pi/512
   cos[431]  =  16'b1100_0111_1011_1110;     //431pi/512
   sin[432]  =  16'b1110_0001_1101_0101;     //432pi/512
   cos[432]  =  16'b1100_0111_1000_1111;     //432pi/512
   sin[433]  =  16'b1110_0010_0010_1101;     //433pi/512
   cos[433]  =  16'b1100_0111_0101_1111;     //433pi/512
   sin[434]  =  16'b1110_0010_1000_0111;     //434pi/512
   cos[434]  =  16'b1100_0111_0011_0001;     //434pi/512
   sin[435]  =  16'b1110_0010_1110_0000;     //435pi/512
   cos[435]  =  16'b1100_0111_0000_0011;     //435pi/512
   sin[436]  =  16'b1110_0011_0011_1010;     //436pi/512
   cos[436]  =  16'b1100_0110_1101_0101;     //436pi/512
   sin[437]  =  16'b1110_0011_1001_0100;     //437pi/512
   cos[437]  =  16'b1100_0110_1010_1000;     //437pi/512
   sin[438]  =  16'b1110_0011_1110_1110;     //438pi/512
   cos[438]  =  16'b1100_0110_0111_1100;     //438pi/512
   sin[439]  =  16'b1110_0100_0100_1000;     //439pi/512
   cos[439]  =  16'b1100_0110_0101_0000;     //439pi/512
   sin[440]  =  16'b1110_0100_1010_0011;     //440pi/512
   cos[440]  =  16'b1100_0110_0010_0101;     //440pi/512
   sin[441]  =  16'b1110_0100_1111_1110;     //441pi/512
   cos[441]  =  16'b1100_0101_1111_1010;     //441pi/512
   sin[442]  =  16'b1110_0101_0101_1001;     //442pi/512
   cos[442]  =  16'b1100_0101_1101_0000;     //442pi/512
   sin[443]  =  16'b1110_0101_1011_0101;     //443pi/512
   cos[443]  =  16'b1100_0101_1010_0111;     //443pi/512
   sin[444]  =  16'b1110_0110_0001_0001;     //444pi/512
   cos[444]  =  16'b1100_0101_0111_1110;     //444pi/512
   sin[445]  =  16'b1110_0110_0110_1101;     //445pi/512
   cos[445]  =  16'b1100_0101_0101_0101;     //445pi/512
   sin[446]  =  16'b1110_0110_1100_1001;     //446pi/512
   cos[446]  =  16'b1100_0101_0010_1101;     //446pi/512
   sin[447]  =  16'b1110_0111_0010_0101;     //447pi/512
   cos[447]  =  16'b1100_0101_0000_0110;     //447pi/512
   sin[448]  =  16'b1110_0111_1000_0010;     //448pi/512
   cos[448]  =  16'b1100_0100_1101_1111;     //448pi/512
   sin[449]  =  16'b1110_0111_1101_1111;     //449pi/512
   cos[449]  =  16'b1100_0100_1011_1001;     //449pi/512
   sin[450]  =  16'b1110_1000_0011_1100;     //450pi/512
   cos[450]  =  16'b1100_0100_1001_0011;     //450pi/512
   sin[451]  =  16'b1110_1000_1001_1010;     //451pi/512
   cos[451]  =  16'b1100_0100_0110_1110;     //451pi/512
   sin[452]  =  16'b1110_1000_1111_0111;     //452pi/512
   cos[452]  =  16'b1100_0100_0100_1010;     //452pi/512
   sin[453]  =  16'b1110_1001_0101_0101;     //453pi/512
   cos[453]  =  16'b1100_0100_0010_0110;     //453pi/512
   sin[454]  =  16'b1110_1001_1011_0100;     //454pi/512
   cos[454]  =  16'b1100_0100_0000_0011;     //454pi/512
   sin[455]  =  16'b1110_1010_0001_0010;     //455pi/512
   cos[455]  =  16'b1100_0011_1110_0000;     //455pi/512
   sin[456]  =  16'b1110_1010_0111_0000;     //456pi/512
   cos[456]  =  16'b1100_0011_1011_1110;     //456pi/512
   sin[457]  =  16'b1110_1010_1100_1111;     //457pi/512
   cos[457]  =  16'b1100_0011_1001_1100;     //457pi/512
   sin[458]  =  16'b1110_1011_0010_1110;     //458pi/512
   cos[458]  =  16'b1100_0011_0111_1011;     //458pi/512
   sin[459]  =  16'b1110_1011_1000_1101;     //459pi/512
   cos[459]  =  16'b1100_0011_0101_1011;     //459pi/512
   sin[460]  =  16'b1110_1011_1110_1101;     //460pi/512
   cos[460]  =  16'b1100_0011_0011_1011;     //460pi/512
   sin[461]  =  16'b1110_1100_0100_1100;     //461pi/512
   cos[461]  =  16'b1100_0011_0001_1100;     //461pi/512
   sin[462]  =  16'b1110_1100_1010_1100;     //462pi/512
   cos[462]  =  16'b1100_0010_1111_1101;     //462pi/512
   sin[463]  =  16'b1110_1101_0000_1100;     //463pi/512
   cos[463]  =  16'b1100_0010_1101_1111;     //463pi/512
   sin[464]  =  16'b1110_1101_0110_1100;     //464pi/512
   cos[464]  =  16'b1100_0010_1100_0001;     //464pi/512
   sin[465]  =  16'b1110_1101_1100_1100;     //465pi/512
   cos[465]  =  16'b1100_0010_1010_0101;     //465pi/512
   sin[466]  =  16'b1110_1110_0010_1101;     //466pi/512
   cos[466]  =  16'b1100_0010_1000_1000;     //466pi/512
   sin[467]  =  16'b1110_1110_1000_1101;     //467pi/512
   cos[467]  =  16'b1100_0010_0110_1101;     //467pi/512
   sin[468]  =  16'b1110_1110_1110_1110;     //468pi/512
   cos[468]  =  16'b1100_0010_0101_0001;     //468pi/512
   sin[469]  =  16'b1110_1111_0100_1111;     //469pi/512
   cos[469]  =  16'b1100_0010_0011_0111;     //469pi/512
   sin[470]  =  16'b1110_1111_1011_0000;     //470pi/512
   cos[470]  =  16'b1100_0010_0001_1101;     //470pi/512
   sin[471]  =  16'b1111_0000_0001_0010;     //471pi/512
   cos[471]  =  16'b1100_0010_0000_0100;     //471pi/512
   sin[472]  =  16'b1111_0000_0111_0011;     //472pi/512
   cos[472]  =  16'b1100_0001_1110_1011;     //472pi/512
   sin[473]  =  16'b1111_0000_1101_0101;     //473pi/512
   cos[473]  =  16'b1100_0001_1101_0011;     //473pi/512
   sin[474]  =  16'b1111_0001_0011_0110;     //474pi/512
   cos[474]  =  16'b1100_0001_1011_1011;     //474pi/512
   sin[475]  =  16'b1111_0001_1001_1000;     //475pi/512
   cos[475]  =  16'b1100_0001_1010_0100;     //475pi/512
   sin[476]  =  16'b1111_0001_1111_1010;     //476pi/512
   cos[476]  =  16'b1100_0001_1000_1110;     //476pi/512
   sin[477]  =  16'b1111_0010_0101_1100;     //477pi/512
   cos[477]  =  16'b1100_0001_0111_1000;     //477pi/512
   sin[478]  =  16'b1111_0010_1011_1111;     //478pi/512
   cos[478]  =  16'b1100_0001_0110_0011;     //478pi/512
   sin[479]  =  16'b1111_0011_0010_0001;     //479pi/512
   cos[479]  =  16'b1100_0001_0100_1111;     //479pi/512
   sin[480]  =  16'b1111_0011_1000_0100;     //480pi/512
   cos[480]  =  16'b1100_0001_0011_1011;     //480pi/512
   sin[481]  =  16'b1111_0011_1110_0110;     //481pi/512
   cos[481]  =  16'b1100_0001_0010_1000;     //481pi/512
   sin[482]  =  16'b1111_0100_0100_1001;     //482pi/512
   cos[482]  =  16'b1100_0001_0001_0101;     //482pi/512
   sin[483]  =  16'b1111_0100_1010_1100;     //483pi/512
   cos[483]  =  16'b1100_0001_0000_0011;     //483pi/512
   sin[484]  =  16'b1111_0101_0000_1111;     //484pi/512
   cos[484]  =  16'b1100_0000_1111_0001;     //484pi/512
   sin[485]  =  16'b1111_0101_0111_0010;     //485pi/512
   cos[485]  =  16'b1100_0000_1110_0000;     //485pi/512
   sin[486]  =  16'b1111_0101_1101_0101;     //486pi/512
   cos[486]  =  16'b1100_0000_1101_0000;     //486pi/512
   sin[487]  =  16'b1111_0110_0011_1001;     //487pi/512
   cos[487]  =  16'b1100_0000_1100_0000;     //487pi/512
   sin[488]  =  16'b1111_0110_1001_1100;     //488pi/512
   cos[488]  =  16'b1100_0000_1011_0001;     //488pi/512
   sin[489]  =  16'b1111_0110_1111_1111;     //489pi/512
   cos[489]  =  16'b1100_0000_1010_0011;     //489pi/512
   sin[490]  =  16'b1111_0111_0110_0011;     //490pi/512
   cos[490]  =  16'b1100_0000_1001_0101;     //490pi/512
   sin[491]  =  16'b1111_0111_1100_0111;     //491pi/512
   cos[491]  =  16'b1100_0000_1000_1000;     //491pi/512
   sin[492]  =  16'b1111_1000_0010_1010;     //492pi/512
   cos[492]  =  16'b1100_0000_0111_1011;     //492pi/512
   sin[493]  =  16'b1111_1000_1000_1110;     //493pi/512
   cos[493]  =  16'b1100_0000_0110_1111;     //493pi/512
   sin[494]  =  16'b1111_1000_1111_0010;     //494pi/512
   cos[494]  =  16'b1100_0000_0110_0100;     //494pi/512
   sin[495]  =  16'b1111_1001_0101_0110;     //495pi/512
   cos[495]  =  16'b1100_0000_0101_1001;     //495pi/512
   sin[496]  =  16'b1111_1001_1011_1010;     //496pi/512
   cos[496]  =  16'b1100_0000_0100_1111;     //496pi/512
   sin[497]  =  16'b1111_1010_0001_1110;     //497pi/512
   cos[497]  =  16'b1100_0000_0100_0101;     //497pi/512
   sin[498]  =  16'b1111_1010_1000_0010;     //498pi/512
   cos[498]  =  16'b1100_0000_0011_1100;     //498pi/512
   sin[499]  =  16'b1111_1010_1110_0110;     //499pi/512
   cos[499]  =  16'b1100_0000_0011_0100;     //499pi/512
   sin[500]  =  16'b1111_1011_0100_1011;     //500pi/512
   cos[500]  =  16'b1100_0000_0010_1100;     //500pi/512
   sin[501]  =  16'b1111_1011_1010_1111;     //501pi/512
   cos[501]  =  16'b1100_0000_0010_0101;     //501pi/512
   sin[502]  =  16'b1111_1100_0001_0011;     //502pi/512
   cos[502]  =  16'b1100_0000_0001_1111;     //502pi/512
   sin[503]  =  16'b1111_1100_0111_1000;     //503pi/512
   cos[503]  =  16'b1100_0000_0001_1001;     //503pi/512
   sin[504]  =  16'b1111_1100_1101_1100;     //504pi/512
   cos[504]  =  16'b1100_0000_0001_0100;     //504pi/512
   sin[505]  =  16'b1111_1101_0100_0000;     //505pi/512
   cos[505]  =  16'b1100_0000_0000_1111;     //505pi/512
   sin[506]  =  16'b1111_1101_1010_0101;     //506pi/512
   cos[506]  =  16'b1100_0000_0000_1011;     //506pi/512
   sin[507]  =  16'b1111_1110_0000_1001;     //507pi/512
   cos[507]  =  16'b1100_0000_0000_1000;     //507pi/512
   sin[508]  =  16'b1111_1110_0110_1110;     //508pi/512
   cos[508]  =  16'b1100_0000_0000_0101;     //508pi/512
   sin[509]  =  16'b1111_1110_1101_0010;     //509pi/512
   cos[509]  =  16'b1100_0000_0000_0011;     //509pi/512
   sin[510]  =  16'b1111_1111_0011_0111;     //510pi/512
   cos[510]  =  16'b1100_0000_0000_0001;     //510pi/512
   sin[511]  =  16'b1111_1111_1001_1011;     //511pi/512
   cos[511]  =  16'b1100_0000_0000_0000;     //511pi/512

   m_sin[0]  =  16'b0000_0000_0000_0000;     //0pi/512
   m_cos[0]  =  16'b0100_0000_0000_0000;     //0pi/512
   m_sin[1]  =  16'b1111_1111_1011_0000;     //1pi/512
   m_cos[1]  =  16'b0011_1111_1111_1111;     //1pi/512
   m_sin[2]  =  16'b1111_1111_0101_1111;     //2pi/512
   m_cos[2]  =  16'b0011_1111_1111_1111;     //2pi/512
   m_sin[3]  =  16'b1111_1111_0000_1111;     //3pi/512
   m_cos[3]  =  16'b0011_1111_1111_1110;     //3pi/512
   m_sin[4]  =  16'b1111_1110_1011_1110;     //4pi/512
   m_cos[4]  =  16'b0011_1111_1111_1100;     //4pi/512
   m_sin[5]  =  16'b1111_1110_0110_1110;     //5pi/512
   m_cos[5]  =  16'b0011_1111_1111_1011;     //5pi/512
   m_sin[6]  =  16'b1111_1110_0001_1110;     //6pi/512
   m_cos[6]  =  16'b0011_1111_1111_1000;     //6pi/512
   m_sin[7]  =  16'b1111_1101_1100_1101;     //7pi/512
   m_cos[7]  =  16'b0011_1111_1111_0110;     //7pi/512
   m_sin[8]  =  16'b1111_1101_0111_1101;     //8pi/512
   m_cos[8]  =  16'b0011_1111_1111_0011;     //8pi/512
   m_sin[9]  =  16'b1111_1101_0010_1100;     //9pi/512
   m_cos[9]  =  16'b0011_1111_1111_0000;     //9pi/512
   m_sin[10]  =  16'b1111_1100_1101_1100;     //10pi/512
   m_cos[10]  =  16'b0011_1111_1110_1100;     //10pi/512
   m_sin[11]  =  16'b1111_1100_1000_1100;     //11pi/512
   m_cos[11]  =  16'b0011_1111_1110_1000;     //11pi/512
   m_sin[12]  =  16'b1111_1100_0011_1011;     //12pi/512
   m_cos[12]  =  16'b0011_1111_1110_0011;     //12pi/512
   m_sin[13]  =  16'b1111_1011_1110_1011;     //13pi/512
   m_cos[13]  =  16'b0011_1111_1101_1110;     //13pi/512
   m_sin[14]  =  16'b1111_1011_1001_1011;     //14pi/512
   m_cos[14]  =  16'b0011_1111_1101_1001;     //14pi/512
   m_sin[15]  =  16'b1111_1011_0100_1011;     //15pi/512
   m_cos[15]  =  16'b0011_1111_1101_0011;     //15pi/512
   m_sin[16]  =  16'b1111_1010_1111_1011;     //16pi/512
   m_cos[16]  =  16'b0011_1111_1100_1101;     //16pi/512
   m_sin[17]  =  16'b1111_1010_1010_1010;     //17pi/512
   m_cos[17]  =  16'b0011_1111_1100_0110;     //17pi/512
   m_sin[18]  =  16'b1111_1010_0101_1010;     //18pi/512
   m_cos[18]  =  16'b0011_1111_1100_0000;     //18pi/512
   m_sin[19]  =  16'b1111_1010_0000_1010;     //19pi/512
   m_cos[19]  =  16'b0011_1111_1011_1000;     //19pi/512
   m_sin[20]  =  16'b1111_1001_1011_1010;     //20pi/512
   m_cos[20]  =  16'b0011_1111_1011_0001;     //20pi/512
   m_sin[21]  =  16'b1111_1001_0110_1010;     //21pi/512
   m_cos[21]  =  16'b0011_1111_1010_1001;     //21pi/512
   m_sin[22]  =  16'b1111_1001_0001_1010;     //22pi/512
   m_cos[22]  =  16'b0011_1111_1010_0000;     //22pi/512
   m_sin[23]  =  16'b1111_1000_1100_1010;     //23pi/512
   m_cos[23]  =  16'b0011_1111_1001_0111;     //23pi/512
   m_sin[24]  =  16'b1111_1000_0111_1010;     //24pi/512
   m_cos[24]  =  16'b0011_1111_1000_1110;     //24pi/512
   m_sin[25]  =  16'b1111_1000_0010_1010;     //25pi/512
   m_cos[25]  =  16'b0011_1111_1000_0100;     //25pi/512
   m_sin[26]  =  16'b1111_0111_1101_1011;     //26pi/512
   m_cos[26]  =  16'b0011_1111_0111_1010;     //26pi/512
   m_sin[27]  =  16'b1111_0111_1000_1011;     //27pi/512
   m_cos[27]  =  16'b0011_1111_0111_0000;     //27pi/512
   m_sin[28]  =  16'b1111_0111_0011_1011;     //28pi/512
   m_cos[28]  =  16'b0011_1111_0110_0101;     //28pi/512
   m_sin[29]  =  16'b1111_0110_1110_1100;     //29pi/512
   m_cos[29]  =  16'b0011_1111_0101_1010;     //29pi/512
   m_sin[30]  =  16'b1111_0110_1001_1100;     //30pi/512
   m_cos[30]  =  16'b0011_1111_0100_1110;     //30pi/512
   m_sin[31]  =  16'b1111_0110_0100_1100;     //31pi/512
   m_cos[31]  =  16'b0011_1111_0100_0010;     //31pi/512
   m_sin[32]  =  16'b1111_0101_1111_1101;     //32pi/512
   m_cos[32]  =  16'b0011_1111_0011_0110;     //32pi/512
   m_sin[33]  =  16'b1111_0101_1010_1110;     //33pi/512
   m_cos[33]  =  16'b0011_1111_0010_1001;     //33pi/512
   m_sin[34]  =  16'b1111_0101_0101_1110;     //34pi/512
   m_cos[34]  =  16'b0011_1111_0001_1100;     //34pi/512
   m_sin[35]  =  16'b1111_0101_0000_1111;     //35pi/512
   m_cos[35]  =  16'b0011_1111_0000_1110;     //35pi/512
   m_sin[36]  =  16'b1111_0100_1100_0000;     //36pi/512
   m_cos[36]  =  16'b0011_1111_0000_0000;     //36pi/512
   m_sin[37]  =  16'b1111_0100_0111_0001;     //37pi/512
   m_cos[37]  =  16'b0011_1110_1111_0010;     //37pi/512
   m_sin[38]  =  16'b1111_0100_0010_0010;     //38pi/512
   m_cos[38]  =  16'b0011_1110_1110_0011;     //38pi/512
   m_sin[39]  =  16'b1111_0011_1101_0011;     //39pi/512
   m_cos[39]  =  16'b0011_1110_1101_0100;     //39pi/512
   m_sin[40]  =  16'b1111_0011_1000_0100;     //40pi/512
   m_cos[40]  =  16'b0011_1110_1100_0101;     //40pi/512
   m_sin[41]  =  16'b1111_0011_0011_0101;     //41pi/512
   m_cos[41]  =  16'b0011_1110_1011_0101;     //41pi/512
   m_sin[42]  =  16'b1111_0010_1110_0110;     //42pi/512
   m_cos[42]  =  16'b0011_1110_1010_0101;     //42pi/512
   m_sin[43]  =  16'b1111_0010_1001_0111;     //43pi/512
   m_cos[43]  =  16'b0011_1110_1001_0100;     //43pi/512
   m_sin[44]  =  16'b1111_0010_0100_1001;     //44pi/512
   m_cos[44]  =  16'b0011_1110_1000_0011;     //44pi/512
   m_sin[45]  =  16'b1111_0001_1111_1010;     //45pi/512
   m_cos[45]  =  16'b0011_1110_0111_0001;     //45pi/512
   m_sin[46]  =  16'b1111_0001_1010_1100;     //46pi/512
   m_cos[46]  =  16'b0011_1110_0110_0000;     //46pi/512
   m_sin[47]  =  16'b1111_0001_0101_1101;     //47pi/512
   m_cos[47]  =  16'b0011_1110_0100_1101;     //47pi/512
   m_sin[48]  =  16'b1111_0001_0000_1111;     //48pi/512
   m_cos[48]  =  16'b0011_1110_0011_1011;     //48pi/512
   m_sin[49]  =  16'b1111_0000_1100_0001;     //49pi/512
   m_cos[49]  =  16'b0011_1110_0010_1000;     //49pi/512
   m_sin[50]  =  16'b1111_0000_0111_0011;     //50pi/512
   m_cos[50]  =  16'b0011_1110_0001_0100;     //50pi/512
   m_sin[51]  =  16'b1111_0000_0010_0101;     //51pi/512
   m_cos[51]  =  16'b0011_1110_0000_0001;     //51pi/512
   m_sin[52]  =  16'b1110_1111_1101_0111;     //52pi/512
   m_cos[52]  =  16'b0011_1101_1110_1101;     //52pi/512
   m_sin[53]  =  16'b1110_1111_1000_1001;     //53pi/512
   m_cos[53]  =  16'b0011_1101_1101_1000;     //53pi/512
   m_sin[54]  =  16'b1110_1111_0011_1100;     //54pi/512
   m_cos[54]  =  16'b0011_1101_1100_0011;     //54pi/512
   m_sin[55]  =  16'b1110_1110_1110_1110;     //55pi/512
   m_cos[55]  =  16'b0011_1101_1010_1110;     //55pi/512
   m_sin[56]  =  16'b1110_1110_1010_0001;     //56pi/512
   m_cos[56]  =  16'b0011_1101_1001_1000;     //56pi/512
   m_sin[57]  =  16'b1110_1110_0101_0011;     //57pi/512
   m_cos[57]  =  16'b0011_1101_1000_0010;     //57pi/512
   m_sin[58]  =  16'b1110_1110_0000_0110;     //58pi/512
   m_cos[58]  =  16'b0011_1101_0110_1100;     //58pi/512
   m_sin[59]  =  16'b1110_1101_1011_1001;     //59pi/512
   m_cos[59]  =  16'b0011_1101_0101_0101;     //59pi/512
   m_sin[60]  =  16'b1110_1101_0110_1100;     //60pi/512
   m_cos[60]  =  16'b0011_1101_0011_1110;     //60pi/512
   m_sin[61]  =  16'b1110_1101_0001_1111;     //61pi/512
   m_cos[61]  =  16'b0011_1101_0010_0110;     //61pi/512
   m_sin[62]  =  16'b1110_1100_1101_0010;     //62pi/512
   m_cos[62]  =  16'b0011_1101_0000_1111;     //62pi/512
   m_sin[63]  =  16'b1110_1100_1000_0110;     //63pi/512
   m_cos[63]  =  16'b0011_1100_1111_0110;     //63pi/512
   m_sin[64]  =  16'b1110_1100_0011_1001;     //64pi/512
   m_cos[64]  =  16'b0011_1100_1101_1110;     //64pi/512
   m_sin[65]  =  16'b1110_1011_1110_1101;     //65pi/512
   m_cos[65]  =  16'b0011_1100_1100_0101;     //65pi/512
   m_sin[66]  =  16'b1110_1011_1010_0000;     //66pi/512
   m_cos[66]  =  16'b0011_1100_1010_1011;     //66pi/512
   m_sin[67]  =  16'b1110_1011_0101_0100;     //67pi/512
   m_cos[67]  =  16'b0011_1100_1001_0001;     //67pi/512
   m_sin[68]  =  16'b1110_1011_0000_1000;     //68pi/512
   m_cos[68]  =  16'b0011_1100_0111_0111;     //68pi/512
   m_sin[69]  =  16'b1110_1010_1011_1100;     //69pi/512
   m_cos[69]  =  16'b0011_1100_0101_1101;     //69pi/512
   m_sin[70]  =  16'b1110_1010_0111_0000;     //70pi/512
   m_cos[70]  =  16'b0011_1100_0100_0010;     //70pi/512
   m_sin[71]  =  16'b1110_1010_0010_0101;     //71pi/512
   m_cos[71]  =  16'b0011_1100_0010_0110;     //71pi/512
   m_sin[72]  =  16'b1110_1001_1101_1001;     //72pi/512
   m_cos[72]  =  16'b0011_1100_0000_1011;     //72pi/512
   m_sin[73]  =  16'b1110_1001_1000_1110;     //73pi/512
   m_cos[73]  =  16'b0011_1011_1110_1111;     //73pi/512
   m_sin[74]  =  16'b1110_1001_0100_0011;     //74pi/512
   m_cos[74]  =  16'b0011_1011_1101_0010;     //74pi/512
   m_sin[75]  =  16'b1110_1000_1111_0111;     //75pi/512
   m_cos[75]  =  16'b0011_1011_1011_0110;     //75pi/512
   m_sin[76]  =  16'b1110_1000_1010_1101;     //76pi/512
   m_cos[76]  =  16'b0011_1011_1001_1001;     //76pi/512
   m_sin[77]  =  16'b1110_1000_0110_0010;     //77pi/512
   m_cos[77]  =  16'b0011_1011_0111_1011;     //77pi/512
   m_sin[78]  =  16'b1110_1000_0001_0111;     //78pi/512
   m_cos[78]  =  16'b0011_1011_0101_1101;     //78pi/512
   m_sin[79]  =  16'b1110_0111_1100_1100;     //79pi/512
   m_cos[79]  =  16'b0011_1011_0011_1111;     //79pi/512
   m_sin[80]  =  16'b1110_0111_1000_0010;     //80pi/512
   m_cos[80]  =  16'b0011_1011_0010_0000;     //80pi/512
   m_sin[81]  =  16'b1110_0111_0011_1000;     //81pi/512
   m_cos[81]  =  16'b0011_1011_0000_0001;     //81pi/512
   m_sin[82]  =  16'b1110_0110_1110_1110;     //82pi/512
   m_cos[82]  =  16'b0011_1010_1110_0010;     //82pi/512
   m_sin[83]  =  16'b1110_0110_1010_0100;     //83pi/512
   m_cos[83]  =  16'b0011_1010_1100_0010;     //83pi/512
   m_sin[84]  =  16'b1110_0110_0101_1010;     //84pi/512
   m_cos[84]  =  16'b0011_1010_1010_0010;     //84pi/512
   m_sin[85]  =  16'b1110_0110_0001_0001;     //85pi/512
   m_cos[85]  =  16'b0011_1010_1000_0010;     //85pi/512
   m_sin[86]  =  16'b1110_0101_1100_0111;     //86pi/512
   m_cos[86]  =  16'b0011_1010_0110_0001;     //86pi/512
   m_sin[87]  =  16'b1110_0101_0111_1110;     //87pi/512
   m_cos[87]  =  16'b0011_1010_0100_0000;     //87pi/512
   m_sin[88]  =  16'b1110_0101_0011_0101;     //88pi/512
   m_cos[88]  =  16'b0011_1010_0001_1111;     //88pi/512
   m_sin[89]  =  16'b1110_0100_1110_1100;     //89pi/512
   m_cos[89]  =  16'b0011_1001_1111_1101;     //89pi/512
   m_sin[90]  =  16'b1110_0100_1010_0011;     //90pi/512
   m_cos[90]  =  16'b0011_1001_1101_1010;     //90pi/512
   m_sin[91]  =  16'b1110_0100_0101_1010;     //91pi/512
   m_cos[91]  =  16'b0011_1001_1011_1000;     //91pi/512
   m_sin[92]  =  16'b1110_0100_0001_0010;     //92pi/512
   m_cos[92]  =  16'b0011_1001_1001_0101;     //92pi/512
   m_sin[93]  =  16'b1110_0011_1100_1010;     //93pi/512
   m_cos[93]  =  16'b0011_1001_0111_0010;     //93pi/512
   m_sin[94]  =  16'b1110_0011_1000_0001;     //94pi/512
   m_cos[94]  =  16'b0011_1001_0100_1110;     //94pi/512
   m_sin[95]  =  16'b1110_0011_0011_1010;     //95pi/512
   m_cos[95]  =  16'b0011_1001_0010_1010;     //95pi/512
   m_sin[96]  =  16'b1110_0010_1111_0010;     //96pi/512
   m_cos[96]  =  16'b0011_1001_0000_0110;     //96pi/512
   m_sin[97]  =  16'b1110_0010_1010_1010;     //97pi/512
   m_cos[97]  =  16'b0011_1000_1110_0001;     //97pi/512
   m_sin[98]  =  16'b1110_0010_0110_0011;     //98pi/512
   m_cos[98]  =  16'b0011_1000_1011_1100;     //98pi/512
   m_sin[99]  =  16'b1110_0010_0001_1100;     //99pi/512
   m_cos[99]  =  16'b0011_1000_1001_0111;     //99pi/512
   m_sin[100]  =  16'b1110_0001_1101_0101;     //100pi/512
   m_cos[100]  =  16'b0011_1000_0111_0001;     //100pi/512
   m_sin[101]  =  16'b1110_0001_1000_1110;     //101pi/512
   m_cos[101]  =  16'b0011_1000_0100_1011;     //101pi/512
   m_sin[102]  =  16'b1110_0001_0100_0111;     //102pi/512
   m_cos[102]  =  16'b0011_1000_0010_0100;     //102pi/512
   m_sin[103]  =  16'b1110_0001_0000_0001;     //103pi/512
   m_cos[103]  =  16'b0011_0111_1111_1110;     //103pi/512
   m_sin[104]  =  16'b1110_0000_1011_1010;     //104pi/512
   m_cos[104]  =  16'b0011_0111_1101_0110;     //104pi/512
   m_sin[105]  =  16'b1110_0000_0111_0100;     //105pi/512
   m_cos[105]  =  16'b0011_0111_1010_1111;     //105pi/512
   m_sin[106]  =  16'b1110_0000_0010_1110;     //106pi/512
   m_cos[106]  =  16'b0011_0111_1000_0111;     //106pi/512
   m_sin[107]  =  16'b1101_1111_1110_1001;     //107pi/512
   m_cos[107]  =  16'b0011_0111_0101_1111;     //107pi/512
   m_sin[108]  =  16'b1101_1111_1010_0011;     //108pi/512
   m_cos[108]  =  16'b0011_0111_0011_0111;     //108pi/512
   m_sin[109]  =  16'b1101_1111_0101_1110;     //109pi/512
   m_cos[109]  =  16'b0011_0111_0000_1110;     //109pi/512
   m_sin[110]  =  16'b1101_1111_0001_1001;     //110pi/512
   m_cos[110]  =  16'b0011_0110_1110_0101;     //110pi/512
   m_sin[111]  =  16'b1101_1110_1101_0100;     //111pi/512
   m_cos[111]  =  16'b0011_0110_1011_1011;     //111pi/512
   m_sin[112]  =  16'b1101_1110_1000_1111;     //112pi/512
   m_cos[112]  =  16'b0011_0110_1001_0001;     //112pi/512
   m_sin[113]  =  16'b1101_1110_0100_1011;     //113pi/512
   m_cos[113]  =  16'b0011_0110_0110_0111;     //113pi/512
   m_sin[114]  =  16'b1101_1110_0000_0111;     //114pi/512
   m_cos[114]  =  16'b0011_0110_0011_1100;     //114pi/512
   m_sin[115]  =  16'b1101_1101_1100_0011;     //115pi/512
   m_cos[115]  =  16'b0011_0110_0001_0010;     //115pi/512
   m_sin[116]  =  16'b1101_1101_0111_1111;     //116pi/512
   m_cos[116]  =  16'b0011_0101_1110_0110;     //116pi/512
   m_sin[117]  =  16'b1101_1101_0011_1011;     //117pi/512
   m_cos[117]  =  16'b0011_0101_1011_1011;     //117pi/512
   m_sin[118]  =  16'b1101_1100_1111_1000;     //118pi/512
   m_cos[118]  =  16'b0011_0101_1000_1111;     //118pi/512
   m_sin[119]  =  16'b1101_1100_1011_0101;     //119pi/512
   m_cos[119]  =  16'b0011_0101_0110_0011;     //119pi/512
   m_sin[120]  =  16'b1101_1100_0111_0010;     //120pi/512
   m_cos[120]  =  16'b0011_0101_0011_0110;     //120pi/512
   m_sin[121]  =  16'b1101_1100_0010_1111;     //121pi/512
   m_cos[121]  =  16'b0011_0101_0000_1001;     //121pi/512
   m_sin[122]  =  16'b1101_1011_1110_1100;     //122pi/512
   m_cos[122]  =  16'b0011_0100_1101_1100;     //122pi/512
   m_sin[123]  =  16'b1101_1011_1010_1010;     //123pi/512
   m_cos[123]  =  16'b0011_0100_1010_1111;     //123pi/512
   m_sin[124]  =  16'b1101_1011_0110_1000;     //124pi/512
   m_cos[124]  =  16'b0011_0100_1000_0001;     //124pi/512
   m_sin[125]  =  16'b1101_1011_0010_0110;     //125pi/512
   m_cos[125]  =  16'b0011_0100_0101_0011;     //125pi/512
   m_sin[126]  =  16'b1101_1010_1110_0100;     //126pi/512
   m_cos[126]  =  16'b0011_0100_0010_0100;     //126pi/512
   m_sin[127]  =  16'b1101_1010_1010_0011;     //127pi/512
   m_cos[127]  =  16'b0011_0011_1111_0110;     //127pi/512
   m_sin[128]  =  16'b1101_1010_0110_0010;     //128pi/512
   m_cos[128]  =  16'b0011_0011_1100_0110;     //128pi/512
   m_sin[129]  =  16'b1101_1010_0010_0001;     //129pi/512
   m_cos[129]  =  16'b0011_0011_1001_0111;     //129pi/512
   m_sin[130]  =  16'b1101_1001_1110_0000;     //130pi/512
   m_cos[130]  =  16'b0011_0011_0110_0111;     //130pi/512
   m_sin[131]  =  16'b1101_1001_1010_0000;     //131pi/512
   m_cos[131]  =  16'b0011_0011_0011_0111;     //131pi/512
   m_sin[132]  =  16'b1101_1001_0101_1111;     //132pi/512
   m_cos[132]  =  16'b0011_0011_0000_0111;     //132pi/512
   m_sin[133]  =  16'b1101_1001_0001_1111;     //133pi/512
   m_cos[133]  =  16'b0011_0010_1101_0110;     //133pi/512
   m_sin[134]  =  16'b1101_1000_1110_0000;     //134pi/512
   m_cos[134]  =  16'b0011_0010_1010_0101;     //134pi/512
   m_sin[135]  =  16'b1101_1000_1010_0000;     //135pi/512
   m_cos[135]  =  16'b0011_0010_0111_0100;     //135pi/512
   m_sin[136]  =  16'b1101_1000_0110_0001;     //136pi/512
   m_cos[136]  =  16'b0011_0010_0100_0010;     //136pi/512
   m_sin[137]  =  16'b1101_1000_0010_0010;     //137pi/512
   m_cos[137]  =  16'b0011_0010_0001_0000;     //137pi/512
   m_sin[138]  =  16'b1101_0111_1110_0011;     //138pi/512
   m_cos[138]  =  16'b0011_0001_1101_1110;     //138pi/512
   m_sin[139]  =  16'b1101_0111_1010_0100;     //139pi/512
   m_cos[139]  =  16'b0011_0001_1010_1011;     //139pi/512
   m_sin[140]  =  16'b1101_0111_0110_0110;     //140pi/512
   m_cos[140]  =  16'b0011_0001_0111_1001;     //140pi/512
   m_sin[141]  =  16'b1101_0111_0010_1000;     //141pi/512
   m_cos[141]  =  16'b0011_0001_0100_0101;     //141pi/512
   m_sin[142]  =  16'b1101_0110_1110_1010;     //142pi/512
   m_cos[142]  =  16'b0011_0001_0001_0010;     //142pi/512
   m_sin[143]  =  16'b1101_0110_1010_1101;     //143pi/512
   m_cos[143]  =  16'b0011_0000_1101_1110;     //143pi/512
   m_sin[144]  =  16'b1101_0110_0110_1111;     //144pi/512
   m_cos[144]  =  16'b0011_0000_1010_1010;     //144pi/512
   m_sin[145]  =  16'b1101_0110_0011_0010;     //145pi/512
   m_cos[145]  =  16'b0011_0000_0111_0110;     //145pi/512
   m_sin[146]  =  16'b1101_0101_1111_0110;     //146pi/512
   m_cos[146]  =  16'b0011_0000_0100_0001;     //146pi/512
   m_sin[147]  =  16'b1101_0101_1011_1001;     //147pi/512
   m_cos[147]  =  16'b0011_0000_0000_1100;     //147pi/512
   m_sin[148]  =  16'b1101_0101_0111_1101;     //148pi/512
   m_cos[148]  =  16'b0010_1111_1101_0111;     //148pi/512
   m_sin[149]  =  16'b1101_0101_0100_0001;     //149pi/512
   m_cos[149]  =  16'b0010_1111_1010_0001;     //149pi/512
   m_sin[150]  =  16'b1101_0101_0000_0101;     //150pi/512
   m_cos[150]  =  16'b0010_1111_0110_1011;     //150pi/512
   m_sin[151]  =  16'b1101_0100_1100_1010;     //151pi/512
   m_cos[151]  =  16'b0010_1111_0011_0101;     //151pi/512
   m_sin[152]  =  16'b1101_0100_1000_1111;     //152pi/512
   m_cos[152]  =  16'b0010_1110_1111_1111;     //152pi/512
   m_sin[153]  =  16'b1101_0100_0101_0100;     //153pi/512
   m_cos[153]  =  16'b0010_1110_1100_1000;     //153pi/512
   m_sin[154]  =  16'b1101_0100_0001_1001;     //154pi/512
   m_cos[154]  =  16'b0010_1110_1001_0001;     //154pi/512
   m_sin[155]  =  16'b1101_0011_1101_1111;     //155pi/512
   m_cos[155]  =  16'b0010_1110_0101_1010;     //155pi/512
   m_sin[156]  =  16'b1101_0011_1010_0100;     //156pi/512
   m_cos[156]  =  16'b0010_1110_0010_0010;     //156pi/512
   m_sin[157]  =  16'b1101_0011_0110_1011;     //157pi/512
   m_cos[157]  =  16'b0010_1101_1110_1010;     //157pi/512
   m_sin[158]  =  16'b1101_0011_0011_0001;     //158pi/512
   m_cos[158]  =  16'b0010_1101_1011_0010;     //158pi/512
   m_sin[159]  =  16'b1101_0010_1111_1000;     //159pi/512
   m_cos[159]  =  16'b0010_1101_0111_1001;     //159pi/512
   m_sin[160]  =  16'b1101_0010_1011_1111;     //160pi/512
   m_cos[160]  =  16'b0010_1101_0100_0001;     //160pi/512
   m_sin[161]  =  16'b1101_0010_1000_0110;     //161pi/512
   m_cos[161]  =  16'b0010_1101_0000_1000;     //161pi/512
   m_sin[162]  =  16'b1101_0010_0100_1110;     //162pi/512
   m_cos[162]  =  16'b0010_1100_1100_1110;     //162pi/512
   m_sin[163]  =  16'b1101_0010_0001_0101;     //163pi/512
   m_cos[163]  =  16'b0010_1100_1001_0101;     //163pi/512
   m_sin[164]  =  16'b1101_0001_1101_1110;     //164pi/512
   m_cos[164]  =  16'b0010_1100_0101_1011;     //164pi/512
   m_sin[165]  =  16'b1101_0001_1010_0110;     //165pi/512
   m_cos[165]  =  16'b0010_1100_0010_0001;     //165pi/512
   m_sin[166]  =  16'b1101_0001_0110_1111;     //166pi/512
   m_cos[166]  =  16'b0010_1011_1110_0111;     //166pi/512
   m_sin[167]  =  16'b1101_0001_0011_1000;     //167pi/512
   m_cos[167]  =  16'b0010_1011_1010_1100;     //167pi/512
   m_sin[168]  =  16'b1101_0001_0000_0001;     //168pi/512
   m_cos[168]  =  16'b0010_1011_0111_0001;     //168pi/512
   m_sin[169]  =  16'b1101_0000_1100_1010;     //169pi/512
   m_cos[169]  =  16'b0010_1011_0011_0110;     //169pi/512
   m_sin[170]  =  16'b1101_0000_1001_0100;     //170pi/512
   m_cos[170]  =  16'b0010_1010_1111_1010;     //170pi/512
   m_sin[171]  =  16'b1101_0000_0101_1110;     //171pi/512
   m_cos[171]  =  16'b0010_1010_1011_1111;     //171pi/512
   m_sin[172]  =  16'b1101_0000_0010_1001;     //172pi/512
   m_cos[172]  =  16'b0010_1010_1000_0011;     //172pi/512
   m_sin[173]  =  16'b1100_1111_1111_0100;     //173pi/512
   m_cos[173]  =  16'b0010_1010_0100_0110;     //173pi/512
   m_sin[174]  =  16'b1100_1111_1011_1111;     //174pi/512
   m_cos[174]  =  16'b0010_1010_0000_1010;     //174pi/512
   m_sin[175]  =  16'b1100_1111_1000_1010;     //175pi/512
   m_cos[175]  =  16'b0010_1001_1100_1101;     //175pi/512
   m_sin[176]  =  16'b1100_1111_0101_0110;     //176pi/512
   m_cos[176]  =  16'b0010_1001_1001_0000;     //176pi/512
   m_sin[177]  =  16'b1100_1111_0010_0001;     //177pi/512
   m_cos[177]  =  16'b0010_1001_0101_0011;     //177pi/512
   m_sin[178]  =  16'b1100_1110_1110_1110;     //178pi/512
   m_cos[178]  =  16'b0010_1001_0001_0101;     //178pi/512
   m_sin[179]  =  16'b1100_1110_1011_1010;     //179pi/512
   m_cos[179]  =  16'b0010_1000_1101_0111;     //179pi/512
   m_sin[180]  =  16'b1100_1110_1000_0111;     //180pi/512
   m_cos[180]  =  16'b0010_1000_1001_1001;     //180pi/512
   m_sin[181]  =  16'b1100_1110_0101_0100;     //181pi/512
   m_cos[181]  =  16'b0010_1000_0101_1011;     //181pi/512
   m_sin[182]  =  16'b1100_1110_0010_0010;     //182pi/512
   m_cos[182]  =  16'b0010_1000_0001_1101;     //182pi/512
   m_sin[183]  =  16'b1100_1101_1110_1111;     //183pi/512
   m_cos[183]  =  16'b0010_0111_1101_1110;     //183pi/512
   m_sin[184]  =  16'b1100_1101_1011_1101;     //184pi/512
   m_cos[184]  =  16'b0010_0111_1001_1111;     //184pi/512
   m_sin[185]  =  16'b1100_1101_1000_1100;     //185pi/512
   m_cos[185]  =  16'b0010_0111_0101_1111;     //185pi/512
   m_sin[186]  =  16'b1100_1101_0101_1010;     //186pi/512
   m_cos[186]  =  16'b0010_0111_0010_0000;     //186pi/512
   m_sin[187]  =  16'b1100_1101_0010_1001;     //187pi/512
   m_cos[187]  =  16'b0010_0110_1110_0000;     //187pi/512
   m_sin[188]  =  16'b1100_1100_1111_1001;     //188pi/512
   m_cos[188]  =  16'b0010_0110_1010_0000;     //188pi/512
   m_sin[189]  =  16'b1100_1100_1100_1000;     //189pi/512
   m_cos[189]  =  16'b0010_0110_0110_0000;     //189pi/512
   m_sin[190]  =  16'b1100_1100_1001_1000;     //190pi/512
   m_cos[190]  =  16'b0010_0110_0001_1111;     //190pi/512
   m_sin[191]  =  16'b1100_1100_0110_1000;     //191pi/512
   m_cos[191]  =  16'b0010_0101_1101_1111;     //191pi/512
   m_sin[192]  =  16'b1100_1100_0011_1001;     //192pi/512
   m_cos[192]  =  16'b0010_0101_1001_1110;     //192pi/512
   m_sin[193]  =  16'b1100_1100_0000_1010;     //193pi/512
   m_cos[193]  =  16'b0010_0101_0101_1101;     //193pi/512
   m_sin[194]  =  16'b1100_1011_1101_1011;     //194pi/512
   m_cos[194]  =  16'b0010_0101_0001_1011;     //194pi/512
   m_sin[195]  =  16'b1100_1011_1010_1101;     //195pi/512
   m_cos[195]  =  16'b0010_0100_1101_1010;     //195pi/512
   m_sin[196]  =  16'b1100_1011_0111_1111;     //196pi/512
   m_cos[196]  =  16'b0010_0100_1001_1000;     //196pi/512
   m_sin[197]  =  16'b1100_1011_0101_0001;     //197pi/512
   m_cos[197]  =  16'b0010_0100_0101_0110;     //197pi/512
   m_sin[198]  =  16'b1100_1011_0010_0011;     //198pi/512
   m_cos[198]  =  16'b0010_0100_0001_0011;     //198pi/512
   m_sin[199]  =  16'b1100_1010_1111_0110;     //199pi/512
   m_cos[199]  =  16'b0010_0011_1101_0001;     //199pi/512
   m_sin[200]  =  16'b1100_1010_1100_1001;     //200pi/512
   m_cos[200]  =  16'b0010_0011_1000_1110;     //200pi/512
   m_sin[201]  =  16'b1100_1010_1001_1101;     //201pi/512
   m_cos[201]  =  16'b0010_0011_0100_1011;     //201pi/512
   m_sin[202]  =  16'b1100_1010_0111_0000;     //202pi/512
   m_cos[202]  =  16'b0010_0011_0000_1000;     //202pi/512
   m_sin[203]  =  16'b1100_1010_0100_0101;     //203pi/512
   m_cos[203]  =  16'b0010_0010_1100_0100;     //203pi/512
   m_sin[204]  =  16'b1100_1010_0001_1001;     //204pi/512
   m_cos[204]  =  16'b0010_0010_1000_0001;     //204pi/512
   m_sin[205]  =  16'b1100_1001_1110_1110;     //205pi/512
   m_cos[205]  =  16'b0010_0010_0011_1101;     //205pi/512
   m_sin[206]  =  16'b1100_1001_1100_0011;     //206pi/512
   m_cos[206]  =  16'b0010_0001_1111_1001;     //206pi/512
   m_sin[207]  =  16'b1100_1001_1001_1001;     //207pi/512
   m_cos[207]  =  16'b0010_0001_1011_0101;     //207pi/512
   m_sin[208]  =  16'b1100_1001_0110_1110;     //208pi/512
   m_cos[208]  =  16'b0010_0001_0111_0000;     //208pi/512
   m_sin[209]  =  16'b1100_1001_0100_0100;     //209pi/512
   m_cos[209]  =  16'b0010_0001_0010_1011;     //209pi/512
   m_sin[210]  =  16'b1100_1001_0001_1011;     //210pi/512
   m_cos[210]  =  16'b0010_0000_1110_0111;     //210pi/512
   m_sin[211]  =  16'b1100_1000_1111_0010;     //211pi/512
   m_cos[211]  =  16'b0010_0000_1010_0001;     //211pi/512
   m_sin[212]  =  16'b1100_1000_1100_1001;     //212pi/512
   m_cos[212]  =  16'b0010_0000_0101_1100;     //212pi/512
   m_sin[213]  =  16'b1100_1000_1010_0000;     //213pi/512
   m_cos[213]  =  16'b0010_0000_0001_0111;     //213pi/512
   m_sin[214]  =  16'b1100_1000_0111_1000;     //214pi/512
   m_cos[214]  =  16'b0001_1111_1101_0001;     //214pi/512
   m_sin[215]  =  16'b1100_1000_0101_0000;     //215pi/512
   m_cos[215]  =  16'b0001_1111_1000_1011;     //215pi/512
   m_sin[216]  =  16'b1100_1000_0010_1001;     //216pi/512
   m_cos[216]  =  16'b0001_1111_0100_0101;     //216pi/512
   m_sin[217]  =  16'b1100_1000_0000_0010;     //217pi/512
   m_cos[217]  =  16'b0001_1110_1111_1111;     //217pi/512
   m_sin[218]  =  16'b1100_0111_1101_1011;     //218pi/512
   m_cos[218]  =  16'b0001_1110_1011_1000;     //218pi/512
   m_sin[219]  =  16'b1100_0111_1011_0101;     //219pi/512
   m_cos[219]  =  16'b0001_1110_0111_0010;     //219pi/512
   m_sin[220]  =  16'b1100_0111_1000_1111;     //220pi/512
   m_cos[220]  =  16'b0001_1110_0010_1011;     //220pi/512
   m_sin[221]  =  16'b1100_0111_0110_1001;     //221pi/512
   m_cos[221]  =  16'b0001_1101_1110_0100;     //221pi/512
   m_sin[222]  =  16'b1100_0111_0100_0011;     //222pi/512
   m_cos[222]  =  16'b0001_1101_1001_1101;     //222pi/512
   m_sin[223]  =  16'b1100_0111_0001_1110;     //223pi/512
   m_cos[223]  =  16'b0001_1101_0101_0101;     //223pi/512
   m_sin[224]  =  16'b1100_0110_1111_1010;     //224pi/512
   m_cos[224]  =  16'b0001_1101_0000_1110;     //224pi/512
   m_sin[225]  =  16'b1100_0110_1101_0101;     //225pi/512
   m_cos[225]  =  16'b0001_1100_1100_0110;     //225pi/512
   m_sin[226]  =  16'b1100_0110_1011_0001;     //226pi/512
   m_cos[226]  =  16'b0001_1100_0111_1110;     //226pi/512
   m_sin[227]  =  16'b1100_0110_1000_1110;     //227pi/512
   m_cos[227]  =  16'b0001_1100_0011_0110;     //227pi/512
   m_sin[228]  =  16'b1100_0110_0110_1011;     //228pi/512
   m_cos[228]  =  16'b0001_1011_1110_1110;     //228pi/512
   m_sin[229]  =  16'b1100_0110_0100_1000;     //229pi/512
   m_cos[229]  =  16'b0001_1011_1010_0101;     //229pi/512
   m_sin[230]  =  16'b1100_0110_0010_0101;     //230pi/512
   m_cos[230]  =  16'b0001_1011_0101_1101;     //230pi/512
   m_sin[231]  =  16'b1100_0110_0000_0011;     //231pi/512
   m_cos[231]  =  16'b0001_1011_0001_0100;     //231pi/512
   m_sin[232]  =  16'b1100_0101_1110_0001;     //232pi/512
   m_cos[232]  =  16'b0001_1010_1100_1011;     //232pi/512
   m_sin[233]  =  16'b1100_0101_1011_1111;     //233pi/512
   m_cos[233]  =  16'b0001_1010_1000_0010;     //233pi/512
   m_sin[234]  =  16'b1100_0101_1001_1110;     //234pi/512
   m_cos[234]  =  16'b0001_1010_0011_1000;     //234pi/512
   m_sin[235]  =  16'b1100_0101_0111_1110;     //235pi/512
   m_cos[235]  =  16'b0001_1001_1110_1111;     //235pi/512
   m_sin[236]  =  16'b1100_0101_0101_1101;     //236pi/512
   m_cos[236]  =  16'b0001_1001_1010_0101;     //236pi/512
   m_sin[237]  =  16'b1100_0101_0011_1101;     //237pi/512
   m_cos[237]  =  16'b0001_1001_0101_1100;     //237pi/512
   m_sin[238]  =  16'b1100_0101_0001_1101;     //238pi/512
   m_cos[238]  =  16'b0001_1001_0001_0010;     //238pi/512
   m_sin[239]  =  16'b1100_0100_1111_1110;     //239pi/512
   m_cos[239]  =  16'b0001_1000_1100_1000;     //239pi/512
   m_sin[240]  =  16'b1100_0100_1101_1111;     //240pi/512
   m_cos[240]  =  16'b0001_1000_0111_1101;     //240pi/512
   m_sin[241]  =  16'b1100_0100_1100_0001;     //241pi/512
   m_cos[241]  =  16'b0001_1000_0011_0011;     //241pi/512
   m_sin[242]  =  16'b1100_0100_1010_0010;     //242pi/512
   m_cos[242]  =  16'b0001_0111_1110_1000;     //242pi/512
   m_sin[243]  =  16'b1100_0100_1000_0100;     //243pi/512
   m_cos[243]  =  16'b0001_0111_1001_1110;     //243pi/512
   m_sin[244]  =  16'b1100_0100_0110_0111;     //244pi/512
   m_cos[244]  =  16'b0001_0111_0101_0011;     //244pi/512
   m_sin[245]  =  16'b1100_0100_0100_1010;     //245pi/512
   m_cos[245]  =  16'b0001_0111_0000_1000;     //245pi/512
   m_sin[246]  =  16'b1100_0100_0010_1101;     //246pi/512
   m_cos[246]  =  16'b0001_0110_1011_1101;     //246pi/512
   m_sin[247]  =  16'b1100_0100_0001_0001;     //247pi/512
   m_cos[247]  =  16'b0001_0110_0111_0010;     //247pi/512
   m_sin[248]  =  16'b1100_0011_1111_0101;     //248pi/512
   m_cos[248]  =  16'b0001_0110_0010_0110;     //248pi/512
   m_sin[249]  =  16'b1100_0011_1101_1001;     //249pi/512
   m_cos[249]  =  16'b0001_0101_1101_1011;     //249pi/512
   m_sin[250]  =  16'b1100_0011_1011_1110;     //250pi/512
   m_cos[250]  =  16'b0001_0101_1000_1111;     //250pi/512
   m_sin[251]  =  16'b1100_0011_1010_0011;     //251pi/512
   m_cos[251]  =  16'b0001_0101_0100_0011;     //251pi/512
   m_sin[252]  =  16'b1100_0011_1000_1000;     //252pi/512
   m_cos[252]  =  16'b0001_0100_1111_0111;     //252pi/512
   m_sin[253]  =  16'b1100_0011_0110_1110;     //253pi/512
   m_cos[253]  =  16'b0001_0100_1010_1011;     //253pi/512
   m_sin[254]  =  16'b1100_0011_0101_0100;     //254pi/512
   m_cos[254]  =  16'b0001_0100_0101_1111;     //254pi/512
   m_sin[255]  =  16'b1100_0011_0011_1011;     //255pi/512
   m_cos[255]  =  16'b0001_0100_0001_0011;     //255pi/512
   m_sin[256]  =  16'b1100_0011_0010_0010;     //256pi/512
   m_cos[256]  =  16'b0001_0011_1100_0110;     //256pi/512
   m_sin[257]  =  16'b1100_0011_0000_1001;     //257pi/512
   m_cos[257]  =  16'b0001_0011_0111_1010;     //257pi/512
   m_sin[258]  =  16'b1100_0010_1111_0001;     //258pi/512
   m_cos[258]  =  16'b0001_0011_0010_1101;     //258pi/512
   m_sin[259]  =  16'b1100_0010_1101_1001;     //259pi/512
   m_cos[259]  =  16'b0001_0010_1110_0000;     //259pi/512
   m_sin[260]  =  16'b1100_0010_1100_0001;     //260pi/512
   m_cos[260]  =  16'b0001_0010_1001_0100;     //260pi/512
   m_sin[261]  =  16'b1100_0010_1010_1010;     //261pi/512
   m_cos[261]  =  16'b0001_0010_0100_0111;     //261pi/512
   m_sin[262]  =  16'b1100_0010_1001_0100;     //262pi/512
   m_cos[262]  =  16'b0001_0001_1111_1001;     //262pi/512
   m_sin[263]  =  16'b1100_0010_0111_1101;     //263pi/512
   m_cos[263]  =  16'b0001_0001_1010_1100;     //263pi/512
   m_sin[264]  =  16'b1100_0010_0110_0111;     //264pi/512
   m_cos[264]  =  16'b0001_0001_0101_1111;     //264pi/512
   m_sin[265]  =  16'b1100_0010_0101_0001;     //265pi/512
   m_cos[265]  =  16'b0001_0001_0001_0001;     //265pi/512
   m_sin[266]  =  16'b1100_0010_0011_1100;     //266pi/512
   m_cos[266]  =  16'b0001_0000_1100_0100;     //266pi/512
   m_sin[267]  =  16'b1100_0010_0010_0111;     //267pi/512
   m_cos[267]  =  16'b0001_0000_0111_0110;     //267pi/512
   m_sin[268]  =  16'b1100_0010_0001_0011;     //268pi/512
   m_cos[268]  =  16'b0001_0000_0010_1000;     //268pi/512
   m_sin[269]  =  16'b1100_0001_1111_1111;     //269pi/512
   m_cos[269]  =  16'b0000_1111_1101_1010;     //269pi/512
   m_sin[270]  =  16'b1100_0001_1110_1011;     //270pi/512
   m_cos[270]  =  16'b0000_1111_1000_1100;     //270pi/512
   m_sin[271]  =  16'b1100_0001_1101_1000;     //271pi/512
   m_cos[271]  =  16'b0000_1111_0011_1110;     //271pi/512
   m_sin[272]  =  16'b1100_0001_1100_0101;     //272pi/512
   m_cos[272]  =  16'b0000_1110_1111_0000;     //272pi/512
   m_sin[273]  =  16'b1100_0001_1011_0010;     //273pi/512
   m_cos[273]  =  16'b0000_1110_1010_0010;     //273pi/512
   m_sin[274]  =  16'b1100_0001_1010_0000;     //274pi/512
   m_cos[274]  =  16'b0000_1110_0101_0100;     //274pi/512
   m_sin[275]  =  16'b1100_0001_1000_1110;     //275pi/512
   m_cos[275]  =  16'b0000_1110_0000_0101;     //275pi/512
   m_sin[276]  =  16'b1100_0001_0111_1101;     //276pi/512
   m_cos[276]  =  16'b0000_1101_1011_0111;     //276pi/512
   m_sin[277]  =  16'b1100_0001_0110_1100;     //277pi/512
   m_cos[277]  =  16'b0000_1101_0110_1000;     //277pi/512
   m_sin[278]  =  16'b1100_0001_0101_1011;     //278pi/512
   m_cos[278]  =  16'b0000_1101_0001_1001;     //278pi/512
   m_sin[279]  =  16'b1100_0001_0100_1011;     //279pi/512
   m_cos[279]  =  16'b0000_1100_1100_1011;     //279pi/512
   m_sin[280]  =  16'b1100_0001_0011_1011;     //280pi/512
   m_cos[280]  =  16'b0000_1100_0111_1100;     //280pi/512
   m_sin[281]  =  16'b1100_0001_0010_1011;     //281pi/512
   m_cos[281]  =  16'b0000_1100_0010_1101;     //281pi/512
   m_sin[282]  =  16'b1100_0001_0001_1100;     //282pi/512
   m_cos[282]  =  16'b0000_1011_1101_1110;     //282pi/512
   m_sin[283]  =  16'b1100_0001_0000_1101;     //283pi/512
   m_cos[283]  =  16'b0000_1011_1000_1111;     //283pi/512
   m_sin[284]  =  16'b1100_0000_1111_1111;     //284pi/512
   m_cos[284]  =  16'b0000_1011_0100_0000;     //284pi/512
   m_sin[285]  =  16'b1100_0000_1111_0001;     //285pi/512
   m_cos[285]  =  16'b0000_1010_1111_0001;     //285pi/512
   m_sin[286]  =  16'b1100_0000_1110_0100;     //286pi/512
   m_cos[286]  =  16'b0000_1010_1010_0001;     //286pi/512
   m_sin[287]  =  16'b1100_0000_1101_0110;     //287pi/512
   m_cos[287]  =  16'b0000_1010_0101_0010;     //287pi/512
   m_sin[288]  =  16'b1100_0000_1100_1010;     //288pi/512
   m_cos[288]  =  16'b0000_1010_0000_0011;     //288pi/512
   m_sin[289]  =  16'b1100_0000_1011_1101;     //289pi/512
   m_cos[289]  =  16'b0000_1001_1011_0011;     //289pi/512
   m_sin[290]  =  16'b1100_0000_1011_0001;     //290pi/512
   m_cos[290]  =  16'b0000_1001_0110_0100;     //290pi/512
   m_sin[291]  =  16'b1100_0000_1010_0110;     //291pi/512
   m_cos[291]  =  16'b0000_1001_0001_0100;     //291pi/512
   m_sin[292]  =  16'b1100_0000_1001_1011;     //292pi/512
   m_cos[292]  =  16'b0000_1000_1100_0100;     //292pi/512
   m_sin[293]  =  16'b1100_0000_1001_0000;     //293pi/512
   m_cos[293]  =  16'b0000_1000_0111_0101;     //293pi/512
   m_sin[294]  =  16'b1100_0000_1000_0101;     //294pi/512
   m_cos[294]  =  16'b0000_1000_0010_0101;     //294pi/512
   m_sin[295]  =  16'b1100_0000_0111_1011;     //295pi/512
   m_cos[295]  =  16'b0000_0111_1101_0101;     //295pi/512
   m_sin[296]  =  16'b1100_0000_0111_0010;     //296pi/512
   m_cos[296]  =  16'b0000_0111_1000_0101;     //296pi/512
   m_sin[297]  =  16'b1100_0000_0110_1000;     //297pi/512
   m_cos[297]  =  16'b0000_0111_0011_0101;     //297pi/512
   m_sin[298]  =  16'b1100_0000_0101_1111;     //298pi/512
   m_cos[298]  =  16'b0000_0110_1110_0101;     //298pi/512
   m_sin[299]  =  16'b1100_0000_0101_0111;     //299pi/512
   m_cos[299]  =  16'b0000_0110_1001_0101;     //299pi/512
   m_sin[300]  =  16'b1100_0000_0100_1111;     //300pi/512
   m_cos[300]  =  16'b0000_0110_0100_0101;     //300pi/512
   m_sin[301]  =  16'b1100_0000_0100_0111;     //301pi/512
   m_cos[301]  =  16'b0000_0101_1111_0101;     //301pi/512
   m_sin[302]  =  16'b1100_0000_0100_0000;     //302pi/512
   m_cos[302]  =  16'b0000_0101_1010_0101;     //302pi/512
   m_sin[303]  =  16'b1100_0000_0011_1001;     //303pi/512
   m_cos[303]  =  16'b0000_0101_0101_0101;     //303pi/512
   m_sin[304]  =  16'b1100_0000_0011_0011;     //304pi/512
   m_cos[304]  =  16'b0000_0101_0000_0101;     //304pi/512
   m_sin[305]  =  16'b1100_0000_0010_1100;     //305pi/512
   m_cos[305]  =  16'b0000_0100_1011_0101;     //305pi/512
   m_sin[306]  =  16'b1100_0000_0010_0111;     //306pi/512
   m_cos[306]  =  16'b0000_0100_0110_0101;     //306pi/512
   m_sin[307]  =  16'b1100_0000_0010_0001;     //307pi/512
   m_cos[307]  =  16'b0000_0100_0001_0100;     //307pi/512
   m_sin[308]  =  16'b1100_0000_0001_1100;     //308pi/512
   m_cos[308]  =  16'b0000_0011_1100_0100;     //308pi/512
   m_sin[309]  =  16'b1100_0000_0001_1000;     //309pi/512
   m_cos[309]  =  16'b0000_0011_0111_0100;     //309pi/512
   m_sin[310]  =  16'b1100_0000_0001_0100;     //310pi/512
   m_cos[310]  =  16'b0000_0011_0010_0011;     //310pi/512
   m_sin[311]  =  16'b1100_0000_0001_0000;     //311pi/512
   m_cos[311]  =  16'b0000_0010_1101_0011;     //311pi/512
   m_sin[312]  =  16'b1100_0000_0000_1101;     //312pi/512
   m_cos[312]  =  16'b0000_0010_1000_0011;     //312pi/512
   m_sin[313]  =  16'b1100_0000_0000_1010;     //313pi/512
   m_cos[313]  =  16'b0000_0010_0011_0010;     //313pi/512
   m_sin[314]  =  16'b1100_0000_0000_0111;     //314pi/512
   m_cos[314]  =  16'b0000_0001_1110_0010;     //314pi/512
   m_sin[315]  =  16'b1100_0000_0000_0101;     //315pi/512
   m_cos[315]  =  16'b0000_0001_1001_0010;     //315pi/512
   m_sin[316]  =  16'b1100_0000_0000_0011;     //316pi/512
   m_cos[316]  =  16'b0000_0001_0100_0001;     //316pi/512
   m_sin[317]  =  16'b1100_0000_0000_0010;     //317pi/512
   m_cos[317]  =  16'b0000_0000_1111_0001;     //317pi/512
   m_sin[318]  =  16'b1100_0000_0000_0001;     //318pi/512
   m_cos[318]  =  16'b0000_0000_1010_0000;     //318pi/512
   m_sin[319]  =  16'b1100_0000_0000_0000;     //319pi/512
   m_cos[319]  =  16'b0000_0000_0101_0000;     //319pi/512
   m_sin[320]  =  16'b1100_0000_0000_0000;     //320pi/512
   m_cos[320]  =  16'b0000_0000_0000_0000;     //320pi/512
   m_sin[321]  =  16'b1100_0000_0000_0000;     //321pi/512
   m_cos[321]  =  16'b1111_1111_1011_0000;     //321pi/512
   m_sin[322]  =  16'b1100_0000_0000_0001;     //322pi/512
   m_cos[322]  =  16'b1111_1111_0101_1111;     //322pi/512
   m_sin[323]  =  16'b1100_0000_0000_0010;     //323pi/512
   m_cos[323]  =  16'b1111_1111_0000_1111;     //323pi/512
   m_sin[324]  =  16'b1100_0000_0000_0011;     //324pi/512
   m_cos[324]  =  16'b1111_1110_1011_1110;     //324pi/512
   m_sin[325]  =  16'b1100_0000_0000_0101;     //325pi/512
   m_cos[325]  =  16'b1111_1110_0110_1110;     //325pi/512
   m_sin[326]  =  16'b1100_0000_0000_0111;     //326pi/512
   m_cos[326]  =  16'b1111_1110_0001_1110;     //326pi/512
   m_sin[327]  =  16'b1100_0000_0000_1010;     //327pi/512
   m_cos[327]  =  16'b1111_1101_1100_1101;     //327pi/512
   m_sin[328]  =  16'b1100_0000_0000_1101;     //328pi/512
   m_cos[328]  =  16'b1111_1101_0111_1101;     //328pi/512
   m_sin[329]  =  16'b1100_0000_0001_0000;     //329pi/512
   m_cos[329]  =  16'b1111_1101_0010_1100;     //329pi/512
   m_sin[330]  =  16'b1100_0000_0001_0100;     //330pi/512
   m_cos[330]  =  16'b1111_1100_1101_1100;     //330pi/512
   m_sin[331]  =  16'b1100_0000_0001_1000;     //331pi/512
   m_cos[331]  =  16'b1111_1100_1000_1100;     //331pi/512
   m_sin[332]  =  16'b1100_0000_0001_1100;     //332pi/512
   m_cos[332]  =  16'b1111_1100_0011_1011;     //332pi/512
   m_sin[333]  =  16'b1100_0000_0010_0001;     //333pi/512
   m_cos[333]  =  16'b1111_1011_1110_1011;     //333pi/512
   m_sin[334]  =  16'b1100_0000_0010_0111;     //334pi/512
   m_cos[334]  =  16'b1111_1011_1001_1011;     //334pi/512
   m_sin[335]  =  16'b1100_0000_0010_1100;     //335pi/512
   m_cos[335]  =  16'b1111_1011_0100_1011;     //335pi/512
   m_sin[336]  =  16'b1100_0000_0011_0011;     //336pi/512
   m_cos[336]  =  16'b1111_1010_1111_1011;     //336pi/512
   m_sin[337]  =  16'b1100_0000_0011_1001;     //337pi/512
   m_cos[337]  =  16'b1111_1010_1010_1010;     //337pi/512
   m_sin[338]  =  16'b1100_0000_0100_0000;     //338pi/512
   m_cos[338]  =  16'b1111_1010_0101_1010;     //338pi/512
   m_sin[339]  =  16'b1100_0000_0100_0111;     //339pi/512
   m_cos[339]  =  16'b1111_1010_0000_1010;     //339pi/512
   m_sin[340]  =  16'b1100_0000_0100_1111;     //340pi/512
   m_cos[340]  =  16'b1111_1001_1011_1010;     //340pi/512
   m_sin[341]  =  16'b1100_0000_0101_0111;     //341pi/512
   m_cos[341]  =  16'b1111_1001_0110_1010;     //341pi/512
   m_sin[342]  =  16'b1100_0000_0101_1111;     //342pi/512
   m_cos[342]  =  16'b1111_1001_0001_1010;     //342pi/512
   m_sin[343]  =  16'b1100_0000_0110_1000;     //343pi/512
   m_cos[343]  =  16'b1111_1000_1100_1010;     //343pi/512
   m_sin[344]  =  16'b1100_0000_0111_0010;     //344pi/512
   m_cos[344]  =  16'b1111_1000_0111_1010;     //344pi/512
   m_sin[345]  =  16'b1100_0000_0111_1011;     //345pi/512
   m_cos[345]  =  16'b1111_1000_0010_1010;     //345pi/512
   m_sin[346]  =  16'b1100_0000_1000_0101;     //346pi/512
   m_cos[346]  =  16'b1111_0111_1101_1011;     //346pi/512
   m_sin[347]  =  16'b1100_0000_1001_0000;     //347pi/512
   m_cos[347]  =  16'b1111_0111_1000_1011;     //347pi/512
   m_sin[348]  =  16'b1100_0000_1001_1011;     //348pi/512
   m_cos[348]  =  16'b1111_0111_0011_1011;     //348pi/512
   m_sin[349]  =  16'b1100_0000_1010_0110;     //349pi/512
   m_cos[349]  =  16'b1111_0110_1110_1100;     //349pi/512
   m_sin[350]  =  16'b1100_0000_1011_0001;     //350pi/512
   m_cos[350]  =  16'b1111_0110_1001_1100;     //350pi/512
   m_sin[351]  =  16'b1100_0000_1011_1101;     //351pi/512
   m_cos[351]  =  16'b1111_0110_0100_1100;     //351pi/512
   m_sin[352]  =  16'b1100_0000_1100_1010;     //352pi/512
   m_cos[352]  =  16'b1111_0101_1111_1101;     //352pi/512
   m_sin[353]  =  16'b1100_0000_1101_0110;     //353pi/512
   m_cos[353]  =  16'b1111_0101_1010_1110;     //353pi/512
   m_sin[354]  =  16'b1100_0000_1110_0100;     //354pi/512
   m_cos[354]  =  16'b1111_0101_0101_1110;     //354pi/512
   m_sin[355]  =  16'b1100_0000_1111_0001;     //355pi/512
   m_cos[355]  =  16'b1111_0101_0000_1111;     //355pi/512
   m_sin[356]  =  16'b1100_0000_1111_1111;     //356pi/512
   m_cos[356]  =  16'b1111_0100_1100_0000;     //356pi/512
   m_sin[357]  =  16'b1100_0001_0000_1101;     //357pi/512
   m_cos[357]  =  16'b1111_0100_0111_0001;     //357pi/512
   m_sin[358]  =  16'b1100_0001_0001_1100;     //358pi/512
   m_cos[358]  =  16'b1111_0100_0010_0010;     //358pi/512
   m_sin[359]  =  16'b1100_0001_0010_1011;     //359pi/512
   m_cos[359]  =  16'b1111_0011_1101_0011;     //359pi/512
   m_sin[360]  =  16'b1100_0001_0011_1011;     //360pi/512
   m_cos[360]  =  16'b1111_0011_1000_0100;     //360pi/512
   m_sin[361]  =  16'b1100_0001_0100_1011;     //361pi/512
   m_cos[361]  =  16'b1111_0011_0011_0101;     //361pi/512
   m_sin[362]  =  16'b1100_0001_0101_1011;     //362pi/512
   m_cos[362]  =  16'b1111_0010_1110_0110;     //362pi/512
   m_sin[363]  =  16'b1100_0001_0110_1100;     //363pi/512
   m_cos[363]  =  16'b1111_0010_1001_0111;     //363pi/512
   m_sin[364]  =  16'b1100_0001_0111_1101;     //364pi/512
   m_cos[364]  =  16'b1111_0010_0100_1001;     //364pi/512
   m_sin[365]  =  16'b1100_0001_1000_1110;     //365pi/512
   m_cos[365]  =  16'b1111_0001_1111_1010;     //365pi/512
   m_sin[366]  =  16'b1100_0001_1010_0000;     //366pi/512
   m_cos[366]  =  16'b1111_0001_1010_1100;     //366pi/512
   m_sin[367]  =  16'b1100_0001_1011_0010;     //367pi/512
   m_cos[367]  =  16'b1111_0001_0101_1101;     //367pi/512
   m_sin[368]  =  16'b1100_0001_1100_0101;     //368pi/512
   m_cos[368]  =  16'b1111_0001_0000_1111;     //368pi/512
   m_sin[369]  =  16'b1100_0001_1101_1000;     //369pi/512
   m_cos[369]  =  16'b1111_0000_1100_0001;     //369pi/512
   m_sin[370]  =  16'b1100_0001_1110_1011;     //370pi/512
   m_cos[370]  =  16'b1111_0000_0111_0011;     //370pi/512
   m_sin[371]  =  16'b1100_0001_1111_1111;     //371pi/512
   m_cos[371]  =  16'b1111_0000_0010_0101;     //371pi/512
   m_sin[372]  =  16'b1100_0010_0001_0011;     //372pi/512
   m_cos[372]  =  16'b1110_1111_1101_0111;     //372pi/512
   m_sin[373]  =  16'b1100_0010_0010_0111;     //373pi/512
   m_cos[373]  =  16'b1110_1111_1000_1001;     //373pi/512
   m_sin[374]  =  16'b1100_0010_0011_1100;     //374pi/512
   m_cos[374]  =  16'b1110_1111_0011_1100;     //374pi/512
   m_sin[375]  =  16'b1100_0010_0101_0001;     //375pi/512
   m_cos[375]  =  16'b1110_1110_1110_1110;     //375pi/512
   m_sin[376]  =  16'b1100_0010_0110_0111;     //376pi/512
   m_cos[376]  =  16'b1110_1110_1010_0001;     //376pi/512
   m_sin[377]  =  16'b1100_0010_0111_1101;     //377pi/512
   m_cos[377]  =  16'b1110_1110_0101_0011;     //377pi/512
   m_sin[378]  =  16'b1100_0010_1001_0100;     //378pi/512
   m_cos[378]  =  16'b1110_1110_0000_0110;     //378pi/512
   m_sin[379]  =  16'b1100_0010_1010_1010;     //379pi/512
   m_cos[379]  =  16'b1110_1101_1011_1001;     //379pi/512
   m_sin[380]  =  16'b1100_0010_1100_0001;     //380pi/512
   m_cos[380]  =  16'b1110_1101_0110_1100;     //380pi/512
   m_sin[381]  =  16'b1100_0010_1101_1001;     //381pi/512
   m_cos[381]  =  16'b1110_1101_0001_1111;     //381pi/512
   m_sin[382]  =  16'b1100_0010_1111_0001;     //382pi/512
   m_cos[382]  =  16'b1110_1100_1101_0010;     //382pi/512
   m_sin[383]  =  16'b1100_0011_0000_1001;     //383pi/512
   m_cos[383]  =  16'b1110_1100_1000_0110;     //383pi/512
   m_sin[384]  =  16'b1100_0011_0010_0010;     //384pi/512
   m_cos[384]  =  16'b1110_1100_0011_1001;     //384pi/512
   m_sin[385]  =  16'b1100_0011_0011_1011;     //385pi/512
   m_cos[385]  =  16'b1110_1011_1110_1101;     //385pi/512
   m_sin[386]  =  16'b1100_0011_0101_0100;     //386pi/512
   m_cos[386]  =  16'b1110_1011_1010_0000;     //386pi/512
   m_sin[387]  =  16'b1100_0011_0110_1110;     //387pi/512
   m_cos[387]  =  16'b1110_1011_0101_0100;     //387pi/512
   m_sin[388]  =  16'b1100_0011_1000_1000;     //388pi/512
   m_cos[388]  =  16'b1110_1011_0000_1000;     //388pi/512
   m_sin[389]  =  16'b1100_0011_1010_0011;     //389pi/512
   m_cos[389]  =  16'b1110_1010_1011_1100;     //389pi/512
   m_sin[390]  =  16'b1100_0011_1011_1110;     //390pi/512
   m_cos[390]  =  16'b1110_1010_0111_0000;     //390pi/512
   m_sin[391]  =  16'b1100_0011_1101_1001;     //391pi/512
   m_cos[391]  =  16'b1110_1010_0010_0101;     //391pi/512
   m_sin[392]  =  16'b1100_0011_1111_0101;     //392pi/512
   m_cos[392]  =  16'b1110_1001_1101_1001;     //392pi/512
   m_sin[393]  =  16'b1100_0100_0001_0001;     //393pi/512
   m_cos[393]  =  16'b1110_1001_1000_1110;     //393pi/512
   m_sin[394]  =  16'b1100_0100_0010_1101;     //394pi/512
   m_cos[394]  =  16'b1110_1001_0100_0011;     //394pi/512
   m_sin[395]  =  16'b1100_0100_0100_1010;     //395pi/512
   m_cos[395]  =  16'b1110_1000_1111_0111;     //395pi/512
   m_sin[396]  =  16'b1100_0100_0110_0111;     //396pi/512
   m_cos[396]  =  16'b1110_1000_1010_1101;     //396pi/512
   m_sin[397]  =  16'b1100_0100_1000_0100;     //397pi/512
   m_cos[397]  =  16'b1110_1000_0110_0010;     //397pi/512
   m_sin[398]  =  16'b1100_0100_1010_0010;     //398pi/512
   m_cos[398]  =  16'b1110_1000_0001_0111;     //398pi/512
   m_sin[399]  =  16'b1100_0100_1100_0001;     //399pi/512
   m_cos[399]  =  16'b1110_0111_1100_1100;     //399pi/512
   m_sin[400]  =  16'b1100_0100_1101_1111;     //400pi/512
   m_cos[400]  =  16'b1110_0111_1000_0010;     //400pi/512
   m_sin[401]  =  16'b1100_0100_1111_1110;     //401pi/512
   m_cos[401]  =  16'b1110_0111_0011_1000;     //401pi/512
   m_sin[402]  =  16'b1100_0101_0001_1101;     //402pi/512
   m_cos[402]  =  16'b1110_0110_1110_1110;     //402pi/512
   m_sin[403]  =  16'b1100_0101_0011_1101;     //403pi/512
   m_cos[403]  =  16'b1110_0110_1010_0100;     //403pi/512
   m_sin[404]  =  16'b1100_0101_0101_1101;     //404pi/512
   m_cos[404]  =  16'b1110_0110_0101_1010;     //404pi/512
   m_sin[405]  =  16'b1100_0101_0111_1110;     //405pi/512
   m_cos[405]  =  16'b1110_0110_0001_0001;     //405pi/512
   m_sin[406]  =  16'b1100_0101_1001_1110;     //406pi/512
   m_cos[406]  =  16'b1110_0101_1100_0111;     //406pi/512
   m_sin[407]  =  16'b1100_0101_1011_1111;     //407pi/512
   m_cos[407]  =  16'b1110_0101_0111_1110;     //407pi/512
   m_sin[408]  =  16'b1100_0101_1110_0001;     //408pi/512
   m_cos[408]  =  16'b1110_0101_0011_0101;     //408pi/512
   m_sin[409]  =  16'b1100_0110_0000_0011;     //409pi/512
   m_cos[409]  =  16'b1110_0100_1110_1100;     //409pi/512
   m_sin[410]  =  16'b1100_0110_0010_0101;     //410pi/512
   m_cos[410]  =  16'b1110_0100_1010_0011;     //410pi/512
   m_sin[411]  =  16'b1100_0110_0100_1000;     //411pi/512
   m_cos[411]  =  16'b1110_0100_0101_1010;     //411pi/512
   m_sin[412]  =  16'b1100_0110_0110_1011;     //412pi/512
   m_cos[412]  =  16'b1110_0100_0001_0010;     //412pi/512
   m_sin[413]  =  16'b1100_0110_1000_1110;     //413pi/512
   m_cos[413]  =  16'b1110_0011_1100_1010;     //413pi/512
   m_sin[414]  =  16'b1100_0110_1011_0001;     //414pi/512
   m_cos[414]  =  16'b1110_0011_1000_0001;     //414pi/512
   m_sin[415]  =  16'b1100_0110_1101_0101;     //415pi/512
   m_cos[415]  =  16'b1110_0011_0011_1010;     //415pi/512
   m_sin[416]  =  16'b1100_0110_1111_1010;     //416pi/512
   m_cos[416]  =  16'b1110_0010_1111_0010;     //416pi/512
   m_sin[417]  =  16'b1100_0111_0001_1110;     //417pi/512
   m_cos[417]  =  16'b1110_0010_1010_1010;     //417pi/512
   m_sin[418]  =  16'b1100_0111_0100_0011;     //418pi/512
   m_cos[418]  =  16'b1110_0010_0110_0011;     //418pi/512
   m_sin[419]  =  16'b1100_0111_0110_1001;     //419pi/512
   m_cos[419]  =  16'b1110_0010_0001_1100;     //419pi/512
   m_sin[420]  =  16'b1100_0111_1000_1111;     //420pi/512
   m_cos[420]  =  16'b1110_0001_1101_0101;     //420pi/512
   m_sin[421]  =  16'b1100_0111_1011_0101;     //421pi/512
   m_cos[421]  =  16'b1110_0001_1000_1110;     //421pi/512
   m_sin[422]  =  16'b1100_0111_1101_1011;     //422pi/512
   m_cos[422]  =  16'b1110_0001_0100_0111;     //422pi/512
   m_sin[423]  =  16'b1100_1000_0000_0010;     //423pi/512
   m_cos[423]  =  16'b1110_0001_0000_0001;     //423pi/512
   m_sin[424]  =  16'b1100_1000_0010_1001;     //424pi/512
   m_cos[424]  =  16'b1110_0000_1011_1010;     //424pi/512
   m_sin[425]  =  16'b1100_1000_0101_0000;     //425pi/512
   m_cos[425]  =  16'b1110_0000_0111_0100;     //425pi/512
   m_sin[426]  =  16'b1100_1000_0111_1000;     //426pi/512
   m_cos[426]  =  16'b1110_0000_0010_1110;     //426pi/512
   m_sin[427]  =  16'b1100_1000_1010_0000;     //427pi/512
   m_cos[427]  =  16'b1101_1111_1110_1001;     //427pi/512
   m_sin[428]  =  16'b1100_1000_1100_1001;     //428pi/512
   m_cos[428]  =  16'b1101_1111_1010_0011;     //428pi/512
   m_sin[429]  =  16'b1100_1000_1111_0010;     //429pi/512
   m_cos[429]  =  16'b1101_1111_0101_1110;     //429pi/512
   m_sin[430]  =  16'b1100_1001_0001_1011;     //430pi/512
   m_cos[430]  =  16'b1101_1111_0001_1001;     //430pi/512
   m_sin[431]  =  16'b1100_1001_0100_0100;     //431pi/512
   m_cos[431]  =  16'b1101_1110_1101_0100;     //431pi/512
   m_sin[432]  =  16'b1100_1001_0110_1110;     //432pi/512
   m_cos[432]  =  16'b1101_1110_1000_1111;     //432pi/512
   m_sin[433]  =  16'b1100_1001_1001_1001;     //433pi/512
   m_cos[433]  =  16'b1101_1110_0100_1011;     //433pi/512
   m_sin[434]  =  16'b1100_1001_1100_0011;     //434pi/512
   m_cos[434]  =  16'b1101_1110_0000_0111;     //434pi/512
   m_sin[435]  =  16'b1100_1001_1110_1110;     //435pi/512
   m_cos[435]  =  16'b1101_1101_1100_0011;     //435pi/512
   m_sin[436]  =  16'b1100_1010_0001_1001;     //436pi/512
   m_cos[436]  =  16'b1101_1101_0111_1111;     //436pi/512
   m_sin[437]  =  16'b1100_1010_0100_0101;     //437pi/512
   m_cos[437]  =  16'b1101_1101_0011_1011;     //437pi/512
   m_sin[438]  =  16'b1100_1010_0111_0000;     //438pi/512
   m_cos[438]  =  16'b1101_1100_1111_1000;     //438pi/512
   m_sin[439]  =  16'b1100_1010_1001_1101;     //439pi/512
   m_cos[439]  =  16'b1101_1100_1011_0101;     //439pi/512
   m_sin[440]  =  16'b1100_1010_1100_1001;     //440pi/512
   m_cos[440]  =  16'b1101_1100_0111_0010;     //440pi/512
   m_sin[441]  =  16'b1100_1010_1111_0110;     //441pi/512
   m_cos[441]  =  16'b1101_1100_0010_1111;     //441pi/512
   m_sin[442]  =  16'b1100_1011_0010_0011;     //442pi/512
   m_cos[442]  =  16'b1101_1011_1110_1100;     //442pi/512
   m_sin[443]  =  16'b1100_1011_0101_0001;     //443pi/512
   m_cos[443]  =  16'b1101_1011_1010_1010;     //443pi/512
   m_sin[444]  =  16'b1100_1011_0111_1111;     //444pi/512
   m_cos[444]  =  16'b1101_1011_0110_1000;     //444pi/512
   m_sin[445]  =  16'b1100_1011_1010_1101;     //445pi/512
   m_cos[445]  =  16'b1101_1011_0010_0110;     //445pi/512
   m_sin[446]  =  16'b1100_1011_1101_1011;     //446pi/512
   m_cos[446]  =  16'b1101_1010_1110_0100;     //446pi/512
   m_sin[447]  =  16'b1100_1100_0000_1010;     //447pi/512
   m_cos[447]  =  16'b1101_1010_1010_0011;     //447pi/512
   m_sin[448]  =  16'b1100_1100_0011_1001;     //448pi/512
   m_cos[448]  =  16'b1101_1010_0110_0010;     //448pi/512
   m_sin[449]  =  16'b1100_1100_0110_1000;     //449pi/512
   m_cos[449]  =  16'b1101_1010_0010_0001;     //449pi/512
   m_sin[450]  =  16'b1100_1100_1001_1000;     //450pi/512
   m_cos[450]  =  16'b1101_1001_1110_0000;     //450pi/512
   m_sin[451]  =  16'b1100_1100_1100_1000;     //451pi/512
   m_cos[451]  =  16'b1101_1001_1010_0000;     //451pi/512
   m_sin[452]  =  16'b1100_1100_1111_1001;     //452pi/512
   m_cos[452]  =  16'b1101_1001_0101_1111;     //452pi/512
   m_sin[453]  =  16'b1100_1101_0010_1001;     //453pi/512
   m_cos[453]  =  16'b1101_1001_0001_1111;     //453pi/512
   m_sin[454]  =  16'b1100_1101_0101_1010;     //454pi/512
   m_cos[454]  =  16'b1101_1000_1110_0000;     //454pi/512
   m_sin[455]  =  16'b1100_1101_1000_1100;     //455pi/512
   m_cos[455]  =  16'b1101_1000_1010_0000;     //455pi/512
   m_sin[456]  =  16'b1100_1101_1011_1101;     //456pi/512
   m_cos[456]  =  16'b1101_1000_0110_0001;     //456pi/512
   m_sin[457]  =  16'b1100_1101_1110_1111;     //457pi/512
   m_cos[457]  =  16'b1101_1000_0010_0010;     //457pi/512
   m_sin[458]  =  16'b1100_1110_0010_0010;     //458pi/512
   m_cos[458]  =  16'b1101_0111_1110_0011;     //458pi/512
   m_sin[459]  =  16'b1100_1110_0101_0100;     //459pi/512
   m_cos[459]  =  16'b1101_0111_1010_0100;     //459pi/512
   m_sin[460]  =  16'b1100_1110_1000_0111;     //460pi/512
   m_cos[460]  =  16'b1101_0111_0110_0110;     //460pi/512
   m_sin[461]  =  16'b1100_1110_1011_1010;     //461pi/512
   m_cos[461]  =  16'b1101_0111_0010_1000;     //461pi/512
   m_sin[462]  =  16'b1100_1110_1110_1110;     //462pi/512
   m_cos[462]  =  16'b1101_0110_1110_1010;     //462pi/512
   m_sin[463]  =  16'b1100_1111_0010_0001;     //463pi/512
   m_cos[463]  =  16'b1101_0110_1010_1101;     //463pi/512
   m_sin[464]  =  16'b1100_1111_0101_0110;     //464pi/512
   m_cos[464]  =  16'b1101_0110_0110_1111;     //464pi/512
   m_sin[465]  =  16'b1100_1111_1000_1010;     //465pi/512
   m_cos[465]  =  16'b1101_0110_0011_0010;     //465pi/512
   m_sin[466]  =  16'b1100_1111_1011_1111;     //466pi/512
   m_cos[466]  =  16'b1101_0101_1111_0110;     //466pi/512
   m_sin[467]  =  16'b1100_1111_1111_0100;     //467pi/512
   m_cos[467]  =  16'b1101_0101_1011_1001;     //467pi/512
   m_sin[468]  =  16'b1101_0000_0010_1001;     //468pi/512
   m_cos[468]  =  16'b1101_0101_0111_1101;     //468pi/512
   m_sin[469]  =  16'b1101_0000_0101_1110;     //469pi/512
   m_cos[469]  =  16'b1101_0101_0100_0001;     //469pi/512
   m_sin[470]  =  16'b1101_0000_1001_0100;     //470pi/512
   m_cos[470]  =  16'b1101_0101_0000_0101;     //470pi/512
   m_sin[471]  =  16'b1101_0000_1100_1010;     //471pi/512
   m_cos[471]  =  16'b1101_0100_1100_1010;     //471pi/512
   m_sin[472]  =  16'b1101_0001_0000_0001;     //472pi/512
   m_cos[472]  =  16'b1101_0100_1000_1111;     //472pi/512
   m_sin[473]  =  16'b1101_0001_0011_1000;     //473pi/512
   m_cos[473]  =  16'b1101_0100_0101_0100;     //473pi/512
   m_sin[474]  =  16'b1101_0001_0110_1111;     //474pi/512
   m_cos[474]  =  16'b1101_0100_0001_1001;     //474pi/512
   m_sin[475]  =  16'b1101_0001_1010_0110;     //475pi/512
   m_cos[475]  =  16'b1101_0011_1101_1111;     //475pi/512
   m_sin[476]  =  16'b1101_0001_1101_1110;     //476pi/512
   m_cos[476]  =  16'b1101_0011_1010_0100;     //476pi/512
   m_sin[477]  =  16'b1101_0010_0001_0101;     //477pi/512
   m_cos[477]  =  16'b1101_0011_0110_1011;     //477pi/512
   m_sin[478]  =  16'b1101_0010_0100_1110;     //478pi/512
   m_cos[478]  =  16'b1101_0011_0011_0001;     //478pi/512
   m_sin[479]  =  16'b1101_0010_1000_0110;     //479pi/512
   m_cos[479]  =  16'b1101_0010_1111_1000;     //479pi/512
   m_sin[480]  =  16'b1101_0010_1011_1111;     //480pi/512
   m_cos[480]  =  16'b1101_0010_1011_1111;     //480pi/512
   m_sin[481]  =  16'b1101_0010_1111_1000;     //481pi/512
   m_cos[481]  =  16'b1101_0010_1000_0110;     //481pi/512
   m_sin[482]  =  16'b1101_0011_0011_0001;     //482pi/512
   m_cos[482]  =  16'b1101_0010_0100_1110;     //482pi/512
   m_sin[483]  =  16'b1101_0011_0110_1011;     //483pi/512
   m_cos[483]  =  16'b1101_0010_0001_0101;     //483pi/512
   m_sin[484]  =  16'b1101_0011_1010_0100;     //484pi/512
   m_cos[484]  =  16'b1101_0001_1101_1110;     //484pi/512
   m_sin[485]  =  16'b1101_0011_1101_1111;     //485pi/512
   m_cos[485]  =  16'b1101_0001_1010_0110;     //485pi/512
   m_sin[486]  =  16'b1101_0100_0001_1001;     //486pi/512
   m_cos[486]  =  16'b1101_0001_0110_1111;     //486pi/512
   m_sin[487]  =  16'b1101_0100_0101_0100;     //487pi/512
   m_cos[487]  =  16'b1101_0001_0011_1000;     //487pi/512
   m_sin[488]  =  16'b1101_0100_1000_1111;     //488pi/512
   m_cos[488]  =  16'b1101_0001_0000_0001;     //488pi/512
   m_sin[489]  =  16'b1101_0100_1100_1010;     //489pi/512
   m_cos[489]  =  16'b1101_0000_1100_1010;     //489pi/512
   m_sin[490]  =  16'b1101_0101_0000_0101;     //490pi/512
   m_cos[490]  =  16'b1101_0000_1001_0100;     //490pi/512
   m_sin[491]  =  16'b1101_0101_0100_0001;     //491pi/512
   m_cos[491]  =  16'b1101_0000_0101_1110;     //491pi/512
   m_sin[492]  =  16'b1101_0101_0111_1101;     //492pi/512
   m_cos[492]  =  16'b1101_0000_0010_1001;     //492pi/512
   m_sin[493]  =  16'b1101_0101_1011_1001;     //493pi/512
   m_cos[493]  =  16'b1100_1111_1111_0100;     //493pi/512
   m_sin[494]  =  16'b1101_0101_1111_0110;     //494pi/512
   m_cos[494]  =  16'b1100_1111_1011_1111;     //494pi/512
   m_sin[495]  =  16'b1101_0110_0011_0010;     //495pi/512
   m_cos[495]  =  16'b1100_1111_1000_1010;     //495pi/512
   m_sin[496]  =  16'b1101_0110_0110_1111;     //496pi/512
   m_cos[496]  =  16'b1100_1111_0101_0110;     //496pi/512
   m_sin[497]  =  16'b1101_0110_1010_1101;     //497pi/512
   m_cos[497]  =  16'b1100_1111_0010_0001;     //497pi/512
   m_sin[498]  =  16'b1101_0110_1110_1010;     //498pi/512
   m_cos[498]  =  16'b1100_1110_1110_1110;     //498pi/512
   m_sin[499]  =  16'b1101_0111_0010_1000;     //499pi/512
   m_cos[499]  =  16'b1100_1110_1011_1010;     //499pi/512
   m_sin[500]  =  16'b1101_0111_0110_0110;     //500pi/512
   m_cos[500]  =  16'b1100_1110_1000_0111;     //500pi/512
   m_sin[501]  =  16'b1101_0111_1010_0100;     //501pi/512
   m_cos[501]  =  16'b1100_1110_0101_0100;     //501pi/512
   m_sin[502]  =  16'b1101_0111_1110_0011;     //502pi/512
   m_cos[502]  =  16'b1100_1110_0010_0010;     //502pi/512
   m_sin[503]  =  16'b1101_1000_0010_0010;     //503pi/512
   m_cos[503]  =  16'b1100_1101_1110_1111;     //503pi/512
   m_sin[504]  =  16'b1101_1000_0110_0001;     //504pi/512
   m_cos[504]  =  16'b1100_1101_1011_1101;     //504pi/512
   m_sin[505]  =  16'b1101_1000_1010_0000;     //505pi/512
   m_cos[505]  =  16'b1100_1101_1000_1100;     //505pi/512
   m_sin[506]  =  16'b1101_1000_1110_0000;     //506pi/512
   m_cos[506]  =  16'b1100_1101_0101_1010;     //506pi/512
   m_sin[507]  =  16'b1101_1001_0001_1111;     //507pi/512
   m_cos[507]  =  16'b1100_1101_0010_1001;     //507pi/512
   m_sin[508]  =  16'b1101_1001_0101_1111;     //508pi/512
   m_cos[508]  =  16'b1100_1100_1111_1001;     //508pi/512
   m_sin[509]  =  16'b1101_1001_1010_0000;     //509pi/512
   m_cos[509]  =  16'b1100_1100_1100_1000;     //509pi/512
   m_sin[510]  =  16'b1101_1001_1110_0000;     //510pi/512
   m_cos[510]  =  16'b1100_1100_1001_1000;     //510pi/512
   m_sin[511]  =  16'b1101_1010_0010_0001;     //511pi/512
   m_cos[511]  =  16'b1100_1100_0110_1000;     //511pi/512
end
endmodule