module  TWIDLE_14_bit_STAGE8_2  #(parameter N = 256, SIZE = 8, bit_width_tw = 14) (
    input                               clk,
    input          [SIZE        -2:0]   rd_ptr_angle,
    input                               en, 

    output reg signed [bit_width_tw-1:0]   cos_data,
    output reg signed [bit_width_tw-1:0]   sin_data
 );

reg signed [bit_width_tw-1:0]  cos  [N/2-1:0];
reg signed [bit_width_tw-1:0]  sin  [N/2-1:0];

localparam  coefficient =  $clog2(256/N);

wire [6:0] rd_ptr = rd_ptr_angle << coefficient;

always @(posedge clk) begin
  if (en) begin
    cos_data <= cos [rd_ptr];
    sin_data <= sin [rd_ptr];
  end
end


initial begin
   sin[0]  =  14'b00100101100111;     //0.2pi/256
   cos[0]  =  14'b00110011110001;     //0.2pi/256
   sin[1]  =  14'b00110011110001;     //0.3pi/256
   cos[1]  =  14'b00100101100111;     //0.3pi/256
   sin[2]  =  14'b00101101010000;     //0.25pi/256
   cos[2]  =  14'b00101101010000;     //0.25pi/256
   sin[3]  =  14'b00111001000001;     //0.35pi/256
   cos[3]  =  14'b00011101000011;     //0.35pi/256
   sin[4]  =  14'b00101001100100;     //0.225pi/256
   cos[4]  =  14'b00110000101010;     //0.225pi/256
   sin[5]  =  14'b00110110100100;     //0.325pi/256
   cos[5]  =  14'b00100001011100;     //0.325pi/256
   sin[6]  =  14'b00110000101010;     //0.275pi/256
   cos[6]  =  14'b00101001100100;     //0.275pi/256
   sin[7]  =  14'b00111011001000;     //0.375pi/256
   cos[7]  =  14'b00011000011111;     //0.375pi/256
   sin[8]  =  14'b00100111100111;     //0.2125pi/256
   cos[8]  =  14'b00110010010000;     //0.2125pi/256
   sin[9]  =  14'b00110101001101;     //0.3125pi/256
   cos[9]  =  14'b00100011100011;     //0.3125pi/256
   sin[10]  =  14'b00101110111111;     //0.2625pi/256
   cos[10]  =  14'b00101011011100;     //0.2625pi/256
   sin[11]  =  14'b00111010000111;     //0.3625pi/256
   cos[11]  =  14'b00011010110010;     //0.3625pi/256
   sin[12]  =  14'b00101011011100;     //0.2375pi/256
   cos[12]  =  14'b00101110111111;     //0.2375pi/256
   sin[13]  =  14'b00110111110101;     //0.3375pi/256
   cos[13]  =  14'b00011111010001;     //0.3375pi/256
   sin[14]  =  14'b00110010010000;     //0.2875pi/256
   cos[14]  =  14'b00100111100111;     //0.2875pi/256
   sin[15]  =  14'b00111100000010;     //0.3875pi/256
   cos[15]  =  14'b00010110001001;     //0.3875pi/256
   sin[16]  =  14'b00100110101000;     //0.20625pi/256
   cos[16]  =  14'b00110011000001;     //0.20625pi/256
   sin[17]  =  14'b00110100100000;     //0.30625pi/256
   cos[17]  =  14'b00100100100110;     //0.30625pi/256
   sin[18]  =  14'b00101110001000;     //0.25625pi/256
   cos[18]  =  14'b00101100010110;     //0.25625pi/256
   sin[19]  =  14'b00111001100101;     //0.35625pi/256
   cos[19]  =  14'b00011011111011;     //0.35625pi/256
   sin[20]  =  14'b00101010100000;     //0.23125pi/256
   cos[20]  =  14'b00101111110101;     //0.23125pi/256
   sin[21]  =  14'b00110111001101;     //0.33125pi/256
   cos[21]  =  14'b00100000010111;     //0.33125pi/256
   sin[22]  =  14'b00110001011110;     //0.28125pi/256
   cos[22]  =  14'b00101000100110;     //0.28125pi/256
   sin[23]  =  14'b00111011100110;     //0.38125pi/256
   cos[23]  =  14'b00010111010100;     //0.38125pi/256
   sin[24]  =  14'b00101000100110;     //0.21875pi/256
   cos[24]  =  14'b00110001011110;     //0.21875pi/256
   sin[25]  =  14'b00110101111001;     //0.31875pi/256
   cos[25]  =  14'b00100010100000;     //0.31875pi/256
   sin[26]  =  14'b00101111110101;     //0.26875pi/256
   cos[26]  =  14'b00101010100000;     //0.26875pi/256
   sin[27]  =  14'b00111010101000;     //0.36875pi/256
   cos[27]  =  14'b00011001101001;     //0.36875pi/256
   sin[28]  =  14'b00101100010110;     //0.24375pi/256
   cos[28]  =  14'b00101110001000;     //0.24375pi/256
   sin[29]  =  14'b00111000011100;     //0.34375pi/256
   cos[29]  =  14'b00011110001010;     //0.34375pi/256
   sin[30]  =  14'b00110011000001;     //0.29375pi/256
   cos[30]  =  14'b00100110101000;     //0.29375pi/256
   sin[31]  =  14'b00111100011101;     //0.39375pi/256
   cos[31]  =  14'b00010100111101;     //0.39375pi/256
   sin[32]  =  14'b00100110000111;     //0.20312pi/256
   cos[32]  =  14'b00110011011001;     //0.20312pi/256
   sin[33]  =  14'b00110100001001;     //0.30313pi/256
   cos[33]  =  14'b00100101000110;     //0.30313pi/256
   sin[34]  =  14'b00101101101100;     //0.25312pi/256
   cos[34]  =  14'b00101100110011;     //0.25312pi/256
   sin[35]  =  14'b00111001010011;     //0.35313pi/256
   cos[35]  =  14'b00011100011111;     //0.35313pi/256
   sin[36]  =  14'b00101010000010;     //0.22813pi/256
   cos[36]  =  14'b00110000010000;     //0.22813pi/256
   sin[37]  =  14'b00110110111001;     //0.32812pi/256
   cos[37]  =  14'b00100000111001;     //0.32812pi/256
   sin[38]  =  14'b00110001000100;     //0.27813pi/256
   cos[38]  =  14'b00101001000101;     //0.27813pi/256
   sin[39]  =  14'b00111011010111;     //0.37813pi/256
   cos[39]  =  14'b00010111111010;     //0.37813pi/256
   sin[40]  =  14'b00101000000111;     //0.21563pi/256
   cos[40]  =  14'b00110001110111;     //0.21563pi/256
   sin[41]  =  14'b00110101100011;     //0.31563pi/256
   cos[41]  =  14'b00100011000010;     //0.31563pi/256
   sin[42]  =  14'b00101111011010;     //0.26562pi/256
   cos[42]  =  14'b00101010111110;     //0.26562pi/256
   sin[43]  =  14'b00111010011000;     //0.36563pi/256
   cos[43]  =  14'b00011010001110;     //0.36563pi/256
   sin[44]  =  14'b00101011111001;     //0.24063pi/256
   cos[44]  =  14'b00101110100100;     //0.24063pi/256
   sin[45]  =  14'b00111000001001;     //0.34063pi/256
   cos[45]  =  14'b00011110101110;     //0.34063pi/256
   sin[46]  =  14'b00110010101001;     //0.29063pi/256
   cos[46]  =  14'b00100111001000;     //0.29063pi/256
   sin[47]  =  14'b00111100010000;     //0.39062pi/256
   cos[47]  =  14'b00010101100011;     //0.39062pi/256
   sin[48]  =  14'b00100111001000;     //0.20938pi/256
   cos[48]  =  14'b00110010101001;     //0.20938pi/256
   sin[49]  =  14'b00110100110111;     //0.30938pi/256
   cos[49]  =  14'b00100100000100;     //0.30938pi/256
   sin[50]  =  14'b00101110100100;     //0.25938pi/256
   cos[50]  =  14'b00101011111001;     //0.25938pi/256
   sin[51]  =  14'b00111001110110;     //0.35938pi/256
   cos[51]  =  14'b00011011010111;     //0.35938pi/256
   sin[52]  =  14'b00101010111110;     //0.23438pi/256
   cos[52]  =  14'b00101111011010;     //0.23438pi/256
   sin[53]  =  14'b00110111100001;     //0.33438pi/256
   cos[53]  =  14'b00011111110100;     //0.33438pi/256
   sin[54]  =  14'b00110001110111;     //0.28437pi/256
   cos[54]  =  14'b00101000000111;     //0.28437pi/256
   sin[55]  =  14'b00111011110100;     //0.38438pi/256
   cos[55]  =  14'b00010110101111;     //0.38438pi/256
   sin[56]  =  14'b00101001000101;     //0.22188pi/256
   cos[56]  =  14'b00110001000100;     //0.22188pi/256
   sin[57]  =  14'b00110110001111;     //0.32188pi/256
   cos[57]  =  14'b00100001111110;     //0.32188pi/256
   sin[58]  =  14'b00110000010000;     //0.27188pi/256
   cos[58]  =  14'b00101010000010;     //0.27188pi/256
   sin[59]  =  14'b00111010111000;     //0.37188pi/256
   cos[59]  =  14'b00011001000100;     //0.37188pi/256
   sin[60]  =  14'b00101100110011;     //0.24688pi/256
   cos[60]  =  14'b00101101101100;     //0.24688pi/256
   sin[61]  =  14'b00111000101111;     //0.34688pi/256
   cos[61]  =  14'b00011101100111;     //0.34688pi/256
   sin[62]  =  14'b00110011011001;     //0.29688pi/256
   cos[62]  =  14'b00100110000111;     //0.29688pi/256
   sin[63]  =  14'b00111100101010;     //0.39688pi/256
   cos[63]  =  14'b00010100010111;     //0.39688pi/256
   sin[64]  =  14'b00100101110111;     //0.20156pi/256
   cos[64]  =  14'b00110011100101;     //0.20156pi/256
   sin[65]  =  14'b00110011111101;     //0.30156pi/256
   cos[65]  =  14'b00100101010111;     //0.30156pi/256
   sin[66]  =  14'b00101101011110;     //0.25156pi/256
   cos[66]  =  14'b00101101000010;     //0.25156pi/256
   sin[67]  =  14'b00111001001010;     //0.35156pi/256
   cos[67]  =  14'b00011100110001;     //0.35156pi/256
   sin[68]  =  14'b00101001110011;     //0.22656pi/256
   cos[68]  =  14'b00110000011101;     //0.22656pi/256
   sin[69]  =  14'b00110110101110;     //0.32656pi/256
   cos[69]  =  14'b00100001001010;     //0.32656pi/256
   sin[70]  =  14'b00110000110111;     //0.27656pi/256
   cos[70]  =  14'b00101001010100;     //0.27656pi/256
   sin[71]  =  14'b00111011001111;     //0.37656pi/256
   cos[71]  =  14'b00011000001100;     //0.37656pi/256
   sin[72]  =  14'b00100111110111;     //0.21406pi/256
   cos[72]  =  14'b00110010000100;     //0.21406pi/256
   sin[73]  =  14'b00110101011000;     //0.31406pi/256
   cos[73]  =  14'b00100011010010;     //0.31406pi/256
   sin[74]  =  14'b00101111001101;     //0.26406pi/256
   cos[74]  =  14'b00101011001101;     //0.26406pi/256
   sin[75]  =  14'b00111010010000;     //0.36406pi/256
   cos[75]  =  14'b00011010100000;     //0.36406pi/256
   sin[76]  =  14'b00101011101011;     //0.23906pi/256
   cos[76]  =  14'b00101110110010;     //0.23906pi/256
   sin[77]  =  14'b00110111111111;     //0.33906pi/256
   cos[77]  =  14'b00011110111111;     //0.33906pi/256
   sin[78]  =  14'b00110010011101;     //0.28906pi/256
   cos[78]  =  14'b00100111010111;     //0.28906pi/256
   sin[79]  =  14'b00111100001001;     //0.38906pi/256
   cos[79]  =  14'b00010101110110;     //0.38906pi/256
   sin[80]  =  14'b00100110111000;     //0.20781pi/256
   cos[80]  =  14'b00110010110101;     //0.20781pi/256
   sin[81]  =  14'b00110100101011;     //0.30781pi/256
   cos[81]  =  14'b00100100010101;     //0.30781pi/256
   sin[82]  =  14'b00101110010110;     //0.25781pi/256
   cos[82]  =  14'b00101100001000;     //0.25781pi/256
   sin[83]  =  14'b00111001101110;     //0.35781pi/256
   cos[83]  =  14'b00011011101001;     //0.35781pi/256
   sin[84]  =  14'b00101010101111;     //0.23281pi/256
   cos[84]  =  14'b00101111101000;     //0.23281pi/256
   sin[85]  =  14'b00110111010111;     //0.33281pi/256
   cos[85]  =  14'b00100000000101;     //0.33281pi/256
   sin[86]  =  14'b00110001101010;     //0.28281pi/256
   cos[86]  =  14'b00101000010110;     //0.28281pi/256
   sin[87]  =  14'b00111011101101;     //0.38281pi/256
   cos[87]  =  14'b00010111000010;     //0.38281pi/256
   sin[88]  =  14'b00101000110101;     //0.22031pi/256
   cos[88]  =  14'b00110001010001;     //0.22031pi/256
   sin[89]  =  14'b00110110000100;     //0.32031pi/256
   cos[89]  =  14'b00100010001111;     //0.32031pi/256
   sin[90]  =  14'b00110000000011;     //0.27031pi/256
   cos[90]  =  14'b00101010010001;     //0.27031pi/256
   sin[91]  =  14'b00111010110000;     //0.37031pi/256
   cos[91]  =  14'b00011001010111;     //0.37031pi/256
   sin[92]  =  14'b00101100100101;     //0.24531pi/256
   cos[92]  =  14'b00101101111010;     //0.24531pi/256
   sin[93]  =  14'b00111000100101;     //0.34531pi/256
   cos[93]  =  14'b00011101111001;     //0.34531pi/256
   sin[94]  =  14'b00110011001101;     //0.29531pi/256
   cos[94]  =  14'b00100110011000;     //0.29531pi/256
   sin[95]  =  14'b00111100100100;     //0.39531pi/256
   cos[95]  =  14'b00010100101010;     //0.39531pi/256
   sin[96]  =  14'b00100110011000;     //0.20469pi/256
   cos[96]  =  14'b00110011001101;     //0.20469pi/256
   sin[97]  =  14'b00110100010100;     //0.30469pi/256
   cos[97]  =  14'b00100100110110;     //0.30469pi/256
   sin[98]  =  14'b00101101111010;     //0.25469pi/256
   cos[98]  =  14'b00101100100101;     //0.25469pi/256
   sin[99]  =  14'b00111001011100;     //0.35469pi/256
   cos[99]  =  14'b00011100001101;     //0.35469pi/256
   sin[100]  =  14'b00101010010001;     //0.22969pi/256
   cos[100]  =  14'b00110000000011;     //0.22969pi/256
   sin[101]  =  14'b00110111000011;     //0.32969pi/256
   cos[101]  =  14'b00100000101000;     //0.32969pi/256
   sin[102]  =  14'b00110001010001;     //0.27969pi/256
   cos[102]  =  14'b00101000110101;     //0.27969pi/256
   sin[103]  =  14'b00111011011110;     //0.37969pi/256
   cos[103]  =  14'b00010111100111;     //0.37969pi/256
   sin[104]  =  14'b00101000010110;     //0.21719pi/256
   cos[104]  =  14'b00110001101010;     //0.21719pi/256
   sin[105]  =  14'b00110101101110;     //0.31719pi/256
   cos[105]  =  14'b00100010110001;     //0.31719pi/256
   sin[106]  =  14'b00101111101000;     //0.26719pi/256
   cos[106]  =  14'b00101010101111;     //0.26719pi/256
   sin[107]  =  14'b00111010100000;     //0.36719pi/256
   cos[107]  =  14'b00011001111011;     //0.36719pi/256
   sin[108]  =  14'b00101100001000;     //0.24219pi/256
   cos[108]  =  14'b00101110010110;     //0.24219pi/256
   sin[109]  =  14'b00111000010010;     //0.34219pi/256
   cos[109]  =  14'b00011110011100;     //0.34219pi/256
   sin[110]  =  14'b00110010110101;     //0.29219pi/256
   cos[110]  =  14'b00100110111000;     //0.29219pi/256
   sin[111]  =  14'b00111100010111;     //0.39219pi/256
   cos[111]  =  14'b00010101010000;     //0.39219pi/256
   sin[112]  =  14'b00100111010111;     //0.21094pi/256
   cos[112]  =  14'b00110010011101;     //0.21094pi/256
   sin[113]  =  14'b00110101000010;     //0.31094pi/256
   cos[113]  =  14'b00100011110100;     //0.31094pi/256
   sin[114]  =  14'b00101110110010;     //0.26094pi/256
   cos[114]  =  14'b00101011101011;     //0.26094pi/256
   sin[115]  =  14'b00111001111111;     //0.36094pi/256
   cos[115]  =  14'b00011011000101;     //0.36094pi/256
   sin[116]  =  14'b00101011001101;     //0.23594pi/256
   cos[116]  =  14'b00101111001101;     //0.23594pi/256
   sin[117]  =  14'b00110111101011;     //0.33594pi/256
   cos[117]  =  14'b00011111100010;     //0.33594pi/256
   sin[118]  =  14'b00110010000100;     //0.28594pi/256
   cos[118]  =  14'b00100111110111;     //0.28594pi/256
   sin[119]  =  14'b00111011111011;     //0.38594pi/256
   cos[119]  =  14'b00010110011100;     //0.38594pi/256
   sin[120]  =  14'b00101001010100;     //0.22344pi/256
   cos[120]  =  14'b00110000110111;     //0.22344pi/256
   sin[121]  =  14'b00110110011001;     //0.32344pi/256
   cos[121]  =  14'b00100001101101;     //0.32344pi/256
   sin[122]  =  14'b00110000011101;     //0.27344pi/256
   cos[122]  =  14'b00101001110011;     //0.27344pi/256
   sin[123]  =  14'b00111011000000;     //0.37344pi/256
   cos[123]  =  14'b00011000110010;     //0.37344pi/256
   sin[124]  =  14'b00101101000010;     //0.24844pi/256
   cos[124]  =  14'b00101101011110;     //0.24844pi/256
   sin[125]  =  14'b00111000111000;     //0.34844pi/256
   cos[125]  =  14'b00011101010101;     //0.34844pi/256
   sin[126]  =  14'b00110011100101;     //0.29844pi/256
   cos[126]  =  14'b00100101110111;     //0.29844pi/256
   sin[127]  =  14'b00111100110001;     //0.39844pi/256
   cos[127]  =  14'b00010100000100;     //0.39844pi/256
end

endmodule