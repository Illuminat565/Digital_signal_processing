module  TWIDLE_12_bit  (
    input   [10:0]   rd_ptr_angle,

    output  signed [11:0]   cos_data,
    output  signed [11:0]   sin_data
 );

wire signed [11:0]  cos  [511:0];
wire signed [11:0]  sin  [511:0];

assign cos_data =    cos [rd_ptr_angle];
assign sin_data =    sin [rd_ptr_angle];


   assign sin[0]  =  12'b000000000000;     //0pi/512
  assign cos[0]  =  12'b010000000000;     //0pi/512
  assign sin[1]  =  12'b111111111010;     //1pi/512
  assign cos[1]  =  12'b001111111111;     //1pi/512
  assign sin[2]  =  12'b111111110011;     //2pi/512
  assign cos[2]  =  12'b001111111111;     //2pi/512
  assign sin[3]  =  12'b111111101101;     //3pi/512
  assign cos[3]  =  12'b001111111111;     //3pi/512
  assign sin[4]  =  12'b111111100111;     //4pi/512
  assign cos[4]  =  12'b001111111111;     //4pi/512
  assign sin[5]  =  12'b111111100001;     //5pi/512
  assign cos[5]  =  12'b001111111111;     //5pi/512
  assign sin[6]  =  12'b111111011010;     //6pi/512
  assign cos[6]  =  12'b001111111111;     //6pi/512
  assign sin[7]  =  12'b111111010100;     //7pi/512
  assign cos[7]  =  12'b001111111111;     //7pi/512
  assign sin[8]  =  12'b111111001110;     //8pi/512
  assign cos[8]  =  12'b001111111110;     //8pi/512
  assign sin[9]  =  12'b111111000111;     //9pi/512
  assign cos[9]  =  12'b001111111110;     //9pi/512
  assign sin[10]  =  12'b111111000001;     //10pi/512
  assign cos[10]  =  12'b001111111110;     //10pi/512
  assign sin[11]  =  12'b111110111011;     //11pi/512
  assign cos[11]  =  12'b001111111101;     //11pi/512
  assign sin[12]  =  12'b111110110101;     //12pi/512
  assign cos[12]  =  12'b001111111101;     //12pi/512
  assign sin[13]  =  12'b111110101110;     //13pi/512
  assign cos[13]  =  12'b001111111100;     //13pi/512
  assign sin[14]  =  12'b111110101000;     //14pi/512
  assign cos[14]  =  12'b001111111100;     //14pi/512
  assign sin[15]  =  12'b111110100010;     //15pi/512
  assign cos[15]  =  12'b001111111011;     //15pi/512
  assign sin[16]  =  12'b111110011100;     //16pi/512
  assign cos[16]  =  12'b001111111011;     //16pi/512
  assign sin[17]  =  12'b111110010101;     //17pi/512
  assign cos[17]  =  12'b001111111010;     //17pi/512
  assign sin[18]  =  12'b111110001111;     //18pi/512
  assign cos[18]  =  12'b001111111001;     //18pi/512
  assign sin[19]  =  12'b111110001001;     //19pi/512
  assign cos[19]  =  12'b001111111001;     //19pi/512
  assign sin[20]  =  12'b111110000011;     //20pi/512
  assign cos[20]  =  12'b001111111000;     //20pi/512
  assign sin[21]  =  12'b111101111100;     //21pi/512
  assign cos[21]  =  12'b001111110111;     //21pi/512
  assign sin[22]  =  12'b111101110110;     //22pi/512
  assign cos[22]  =  12'b001111110110;     //22pi/512
  assign sin[23]  =  12'b111101110000;     //23pi/512
  assign cos[23]  =  12'b001111110101;     //23pi/512
  assign sin[24]  =  12'b111101101010;     //24pi/512
  assign cos[24]  =  12'b001111110100;     //24pi/512
  assign sin[25]  =  12'b111101100100;     //25pi/512
  assign cos[25]  =  12'b001111110011;     //25pi/512
  assign sin[26]  =  12'b111101011101;     //26pi/512
  assign cos[26]  =  12'b001111110010;     //26pi/512
  assign sin[27]  =  12'b111101010111;     //27pi/512
  assign cos[27]  =  12'b001111110001;     //27pi/512
  assign sin[28]  =  12'b111101010001;     //28pi/512
  assign cos[28]  =  12'b001111110000;     //28pi/512
  assign sin[29]  =  12'b111101001011;     //29pi/512
  assign cos[29]  =  12'b001111101111;     //29pi/512
  assign sin[30]  =  12'b111101000101;     //30pi/512
  assign cos[30]  =  12'b001111101110;     //30pi/512
  assign sin[31]  =  12'b111100111110;     //31pi/512
  assign cos[31]  =  12'b001111101101;     //31pi/512
  assign sin[32]  =  12'b111100111000;     //32pi/512
  assign cos[32]  =  12'b001111101100;     //32pi/512
  assign sin[33]  =  12'b111100110010;     //33pi/512
  assign cos[33]  =  12'b001111101011;     //33pi/512
  assign sin[34]  =  12'b111100101100;     //34pi/512
  assign cos[34]  =  12'b001111101001;     //34pi/512
  assign sin[35]  =  12'b111100100110;     //35pi/512
  assign cos[35]  =  12'b001111101000;     //35pi/512
  assign sin[36]  =  12'b111100100000;     //36pi/512
  assign cos[36]  =  12'b001111100111;     //36pi/512
  assign sin[37]  =  12'b111100011010;     //37pi/512
  assign cos[37]  =  12'b001111100101;     //37pi/512
  assign sin[38]  =  12'b111100010011;     //38pi/512
  assign cos[38]  =  12'b001111100100;     //38pi/512
  assign sin[39]  =  12'b111100001101;     //39pi/512
  assign cos[39]  =  12'b001111100010;     //39pi/512
  assign sin[40]  =  12'b111100000111;     //40pi/512
  assign cos[40]  =  12'b001111100001;     //40pi/512
  assign sin[41]  =  12'b111100000001;     //41pi/512
  assign cos[41]  =  12'b001111011111;     //41pi/512
  assign sin[42]  =  12'b111011111011;     //42pi/512
  assign cos[42]  =  12'b001111011110;     //42pi/512
  assign sin[43]  =  12'b111011110101;     //43pi/512
  assign cos[43]  =  12'b001111011100;     //43pi/512
  assign sin[44]  =  12'b111011101111;     //44pi/512
  assign cos[44]  =  12'b001111011010;     //44pi/512
  assign sin[45]  =  12'b111011101001;     //45pi/512
  assign cos[45]  =  12'b001111011001;     //45pi/512
  assign sin[46]  =  12'b111011100011;     //46pi/512
  assign cos[46]  =  12'b001111010111;     //46pi/512
  assign sin[47]  =  12'b111011011101;     //47pi/512
  assign cos[47]  =  12'b001111010101;     //47pi/512
  assign sin[48]  =  12'b111011010111;     //48pi/512
  assign cos[48]  =  12'b001111010011;     //48pi/512
  assign sin[49]  =  12'b111011010001;     //49pi/512
  assign cos[49]  =  12'b001111010010;     //49pi/512
  assign sin[50]  =  12'b111011001011;     //50pi/512
  assign cos[50]  =  12'b001111010000;     //50pi/512
  assign sin[51]  =  12'b111011000101;     //51pi/512
  assign cos[51]  =  12'b001111001110;     //51pi/512
  assign sin[52]  =  12'b111010111111;     //52pi/512
  assign cos[52]  =  12'b001111001100;     //52pi/512
  assign sin[53]  =  12'b111010111001;     //53pi/512
  assign cos[53]  =  12'b001111001010;     //53pi/512
  assign sin[54]  =  12'b111010110011;     //54pi/512
  assign cos[54]  =  12'b001111001000;     //54pi/512
  assign sin[55]  =  12'b111010101101;     //55pi/512
  assign cos[55]  =  12'b001111000110;     //55pi/512
  assign sin[56]  =  12'b111010100111;     //56pi/512
  assign cos[56]  =  12'b001111000100;     //56pi/512
  assign sin[57]  =  12'b111010100001;     //57pi/512
  assign cos[57]  =  12'b001111000010;     //57pi/512
  assign sin[58]  =  12'b111010011011;     //58pi/512
  assign cos[58]  =  12'b001110111111;     //58pi/512
  assign sin[59]  =  12'b111010010101;     //59pi/512
  assign cos[59]  =  12'b001110111101;     //59pi/512
  assign sin[60]  =  12'b111010001111;     //60pi/512
  assign cos[60]  =  12'b001110111011;     //60pi/512
  assign sin[61]  =  12'b111010001010;     //61pi/512
  assign cos[61]  =  12'b001110111001;     //61pi/512
  assign sin[62]  =  12'b111010000100;     //62pi/512
  assign cos[62]  =  12'b001110110110;     //62pi/512
  assign sin[63]  =  12'b111001111110;     //63pi/512
  assign cos[63]  =  12'b001110110100;     //63pi/512
  assign sin[64]  =  12'b111001111000;     //64pi/512
  assign cos[64]  =  12'b001110110010;     //64pi/512
  assign sin[65]  =  12'b111001110010;     //65pi/512
  assign cos[65]  =  12'b001110101111;     //65pi/512
  assign sin[66]  =  12'b111001101101;     //66pi/512
  assign cos[66]  =  12'b001110101101;     //66pi/512
  assign sin[67]  =  12'b111001100111;     //67pi/512
  assign cos[67]  =  12'b001110101010;     //67pi/512
  assign sin[68]  =  12'b111001100001;     //68pi/512
  assign cos[68]  =  12'b001110101000;     //68pi/512
  assign sin[69]  =  12'b111001011011;     //69pi/512
  assign cos[69]  =  12'b001110100101;     //69pi/512
  assign sin[70]  =  12'b111001010110;     //70pi/512
  assign cos[70]  =  12'b001110100010;     //70pi/512
  assign sin[71]  =  12'b111001010000;     //71pi/512
  assign cos[71]  =  12'b001110100000;     //71pi/512
  assign sin[72]  =  12'b111001001010;     //72pi/512
  assign cos[72]  =  12'b001110011101;     //72pi/512
  assign sin[73]  =  12'b111001000101;     //73pi/512
  assign cos[73]  =  12'b001110011010;     //73pi/512
  assign sin[74]  =  12'b111000111111;     //74pi/512
  assign cos[74]  =  12'b001110011000;     //74pi/512
  assign sin[75]  =  12'b111000111001;     //75pi/512
  assign cos[75]  =  12'b001110010101;     //75pi/512
  assign sin[76]  =  12'b111000110100;     //76pi/512
  assign cos[76]  =  12'b001110010010;     //76pi/512
  assign sin[77]  =  12'b111000101110;     //77pi/512
  assign cos[77]  =  12'b001110001111;     //77pi/512
  assign sin[78]  =  12'b111000101000;     //78pi/512
  assign cos[78]  =  12'b001110001100;     //78pi/512
  assign sin[79]  =  12'b111000100011;     //79pi/512
  assign cos[79]  =  12'b001110001010;     //79pi/512
  assign sin[80]  =  12'b111000011101;     //80pi/512
  assign cos[80]  =  12'b001110000111;     //80pi/512
  assign sin[81]  =  12'b111000011000;     //81pi/512
  assign cos[81]  =  12'b001110000100;     //81pi/512
  assign sin[82]  =  12'b111000010010;     //82pi/512
  assign cos[82]  =  12'b001110000001;     //82pi/512
  assign sin[83]  =  12'b111000001101;     //83pi/512
  assign cos[83]  =  12'b001101111110;     //83pi/512
  assign sin[84]  =  12'b111000000111;     //84pi/512
  assign cos[84]  =  12'b001101111010;     //84pi/512
  assign sin[85]  =  12'b111000000010;     //85pi/512
  assign cos[85]  =  12'b001101110111;     //85pi/512
  assign sin[86]  =  12'b110111111100;     //86pi/512
  assign cos[86]  =  12'b001101110100;     //86pi/512
  assign sin[87]  =  12'b110111110111;     //87pi/512
  assign cos[87]  =  12'b001101110001;     //87pi/512
  assign sin[88]  =  12'b110111110010;     //88pi/512
  assign cos[88]  =  12'b001101101110;     //88pi/512
  assign sin[89]  =  12'b110111101100;     //89pi/512
  assign cos[89]  =  12'b001101101011;     //89pi/512
  assign sin[90]  =  12'b110111100111;     //90pi/512
  assign cos[90]  =  12'b001101100111;     //90pi/512
  assign sin[91]  =  12'b110111100001;     //91pi/512
  assign cos[91]  =  12'b001101100100;     //91pi/512
  assign sin[92]  =  12'b110111011100;     //92pi/512
  assign cos[92]  =  12'b001101100001;     //92pi/512
  assign sin[93]  =  12'b110111010111;     //93pi/512
  assign cos[93]  =  12'b001101011101;     //93pi/512
  assign sin[94]  =  12'b110111010010;     //94pi/512
  assign cos[94]  =  12'b001101011010;     //94pi/512
  assign sin[95]  =  12'b110111001100;     //95pi/512
  assign cos[95]  =  12'b001101010110;     //95pi/512
  assign sin[96]  =  12'b110111000111;     //96pi/512
  assign cos[96]  =  12'b001101010011;     //96pi/512
  assign sin[97]  =  12'b110111000010;     //97pi/512
  assign cos[97]  =  12'b001101001111;     //97pi/512
  assign sin[98]  =  12'b110110111101;     //98pi/512
  assign cos[98]  =  12'b001101001100;     //98pi/512
  assign sin[99]  =  12'b110110111000;     //99pi/512
  assign cos[99]  =  12'b001101001000;     //99pi/512
  assign sin[100]  =  12'b110110110010;     //100pi/512
  assign cos[100]  =  12'b001101000101;     //100pi/512
  assign sin[101]  =  12'b110110101101;     //101pi/512
  assign cos[101]  =  12'b001101000001;     //101pi/512
  assign sin[102]  =  12'b110110101000;     //102pi/512
  assign cos[102]  =  12'b001100111101;     //102pi/512
  assign sin[103]  =  12'b110110100011;     //103pi/512
  assign cos[103]  =  12'b001100111010;     //103pi/512
  assign sin[104]  =  12'b110110011110;     //104pi/512
  assign cos[104]  =  12'b001100110110;     //104pi/512
  assign sin[105]  =  12'b110110011001;     //105pi/512
  assign cos[105]  =  12'b001100110010;     //105pi/512
  assign sin[106]  =  12'b110110010100;     //106pi/512
  assign cos[106]  =  12'b001100101110;     //106pi/512
  assign sin[107]  =  12'b110110001111;     //107pi/512
  assign cos[107]  =  12'b001100101011;     //107pi/512
  assign sin[108]  =  12'b110110001010;     //108pi/512
  assign cos[108]  =  12'b001100100111;     //108pi/512
  assign sin[109]  =  12'b110110000101;     //109pi/512
  assign cos[109]  =  12'b001100100011;     //109pi/512
  assign sin[110]  =  12'b110110000000;     //110pi/512
  assign cos[110]  =  12'b001100011111;     //110pi/512
  assign sin[111]  =  12'b110101111011;     //111pi/512
  assign cos[111]  =  12'b001100011011;     //111pi/512
  assign sin[112]  =  12'b110101110110;     //112pi/512
  assign cos[112]  =  12'b001100010111;     //112pi/512
  assign sin[113]  =  12'b110101110010;     //113pi/512
  assign cos[113]  =  12'b001100010011;     //113pi/512
  assign sin[114]  =  12'b110101101101;     //114pi/512
  assign cos[114]  =  12'b001100001111;     //114pi/512
  assign sin[115]  =  12'b110101101000;     //115pi/512
  assign cos[115]  =  12'b001100001011;     //115pi/512
  assign sin[116]  =  12'b110101100011;     //116pi/512
  assign cos[116]  =  12'b001100000111;     //116pi/512
  assign sin[117]  =  12'b110101011110;     //117pi/512
  assign cos[117]  =  12'b001100000011;     //117pi/512
  assign sin[118]  =  12'b110101011010;     //118pi/512
  assign cos[118]  =  12'b001011111111;     //118pi/512
  assign sin[119]  =  12'b110101010101;     //119pi/512
  assign cos[119]  =  12'b001011111010;     //119pi/512
  assign sin[120]  =  12'b110101010000;     //120pi/512
  assign cos[120]  =  12'b001011110110;     //120pi/512
  assign sin[121]  =  12'b110101001100;     //121pi/512
  assign cos[121]  =  12'b001011110010;     //121pi/512
  assign sin[122]  =  12'b110101000111;     //122pi/512
  assign cos[122]  =  12'b001011101110;     //122pi/512
  assign sin[123]  =  12'b110101000010;     //123pi/512
  assign cos[123]  =  12'b001011101001;     //123pi/512
  assign sin[124]  =  12'b110100111110;     //124pi/512
  assign cos[124]  =  12'b001011100101;     //124pi/512
  assign sin[125]  =  12'b110100111001;     //125pi/512
  assign cos[125]  =  12'b001011100001;     //125pi/512
  assign sin[126]  =  12'b110100110101;     //126pi/512
  assign cos[126]  =  12'b001011011100;     //126pi/512
  assign sin[127]  =  12'b110100110000;     //127pi/512
  assign cos[127]  =  12'b001011011000;     //127pi/512
  assign sin[128]  =  12'b110100101100;     //128pi/512
  assign cos[128]  =  12'b001011010100;     //128pi/512
  assign sin[129]  =  12'b110100100111;     //129pi/512
  assign cos[129]  =  12'b001011001111;     //129pi/512
  assign sin[130]  =  12'b110100100011;     //130pi/512
  assign cos[130]  =  12'b001011001011;     //130pi/512
  assign sin[131]  =  12'b110100011111;     //131pi/512
  assign cos[131]  =  12'b001011000110;     //131pi/512
  assign sin[132]  =  12'b110100011010;     //132pi/512
  assign cos[132]  =  12'b001011000010;     //132pi/512
  assign sin[133]  =  12'b110100010110;     //133pi/512
  assign cos[133]  =  12'b001010111101;     //133pi/512
  assign sin[134]  =  12'b110100010010;     //134pi/512
  assign cos[134]  =  12'b001010111000;     //134pi/512
  assign sin[135]  =  12'b110100001101;     //135pi/512
  assign cos[135]  =  12'b001010110100;     //135pi/512
  assign sin[136]  =  12'b110100001001;     //136pi/512
  assign cos[136]  =  12'b001010101111;     //136pi/512
  assign sin[137]  =  12'b110100000101;     //137pi/512
  assign cos[137]  =  12'b001010101011;     //137pi/512
  assign sin[138]  =  12'b110100000001;     //138pi/512
  assign cos[138]  =  12'b001010100110;     //138pi/512
  assign sin[139]  =  12'b110011111101;     //139pi/512
  assign cos[139]  =  12'b001010100001;     //139pi/512
  assign sin[140]  =  12'b110011111001;     //140pi/512
  assign cos[140]  =  12'b001010011100;     //140pi/512
  assign sin[141]  =  12'b110011110101;     //141pi/512
  assign cos[141]  =  12'b001010011000;     //141pi/512
  assign sin[142]  =  12'b110011110000;     //142pi/512
  assign cos[142]  =  12'b001010010011;     //142pi/512
  assign sin[143]  =  12'b110011101100;     //143pi/512
  assign cos[143]  =  12'b001010001110;     //143pi/512
  assign sin[144]  =  12'b110011101000;     //144pi/512
  assign cos[144]  =  12'b001010001001;     //144pi/512
  assign sin[145]  =  12'b110011100100;     //145pi/512
  assign cos[145]  =  12'b001010000100;     //145pi/512
  assign sin[146]  =  12'b110011100001;     //146pi/512
  assign cos[146]  =  12'b001001111111;     //146pi/512
  assign sin[147]  =  12'b110011011101;     //147pi/512
  assign cos[147]  =  12'b001001111010;     //147pi/512
  assign sin[148]  =  12'b110011011001;     //148pi/512
  assign cos[148]  =  12'b001001110101;     //148pi/512
  assign sin[149]  =  12'b110011010101;     //149pi/512
  assign cos[149]  =  12'b001001110001;     //149pi/512
  assign sin[150]  =  12'b110011010001;     //150pi/512
  assign cos[150]  =  12'b001001101100;     //150pi/512
  assign sin[151]  =  12'b110011001101;     //151pi/512
  assign cos[151]  =  12'b001001100111;     //151pi/512
  assign sin[152]  =  12'b110011001010;     //152pi/512
  assign cos[152]  =  12'b001001100001;     //152pi/512
  assign sin[153]  =  12'b110011000110;     //153pi/512
  assign cos[153]  =  12'b001001011100;     //153pi/512
  assign sin[154]  =  12'b110011000010;     //154pi/512
  assign cos[154]  =  12'b001001010111;     //154pi/512
  assign sin[155]  =  12'b110010111110;     //155pi/512
  assign cos[155]  =  12'b001001010010;     //155pi/512
  assign sin[156]  =  12'b110010111011;     //156pi/512
  assign cos[156]  =  12'b001001001101;     //156pi/512
  assign sin[157]  =  12'b110010110111;     //157pi/512
  assign cos[157]  =  12'b001001001000;     //157pi/512
  assign sin[158]  =  12'b110010110100;     //158pi/512
  assign cos[158]  =  12'b001001000011;     //158pi/512
  assign sin[159]  =  12'b110010110000;     //159pi/512
  assign cos[159]  =  12'b001000111110;     //159pi/512
  assign sin[160]  =  12'b110010101101;     //160pi/512
  assign cos[160]  =  12'b001000111000;     //160pi/512
  assign sin[161]  =  12'b110010101001;     //161pi/512
  assign cos[161]  =  12'b001000110011;     //161pi/512
  assign sin[162]  =  12'b110010100110;     //162pi/512
  assign cos[162]  =  12'b001000101110;     //162pi/512
  assign sin[163]  =  12'b110010100010;     //163pi/512
  assign cos[163]  =  12'b001000101001;     //163pi/512
  assign sin[164]  =  12'b110010011111;     //164pi/512
  assign cos[164]  =  12'b001000100011;     //164pi/512
  assign sin[165]  =  12'b110010011100;     //165pi/512
  assign cos[165]  =  12'b001000011110;     //165pi/512
  assign sin[166]  =  12'b110010011000;     //166pi/512
  assign cos[166]  =  12'b001000011001;     //166pi/512
  assign sin[167]  =  12'b110010010101;     //167pi/512
  assign cos[167]  =  12'b001000010011;     //167pi/512
  assign sin[168]  =  12'b110010010010;     //168pi/512
  assign cos[168]  =  12'b001000001110;     //168pi/512
  assign sin[169]  =  12'b110010001110;     //169pi/512
  assign cos[169]  =  12'b001000001001;     //169pi/512
  assign sin[170]  =  12'b110010001011;     //170pi/512
  assign cos[170]  =  12'b001000000011;     //170pi/512
  assign sin[171]  =  12'b110010001000;     //171pi/512
  assign cos[171]  =  12'b000111111110;     //171pi/512
  assign sin[172]  =  12'b110010000101;     //172pi/512
  assign cos[172]  =  12'b000111111000;     //172pi/512
  assign sin[173]  =  12'b110010000010;     //173pi/512
  assign cos[173]  =  12'b000111110011;     //173pi/512
  assign sin[174]  =  12'b110001111111;     //174pi/512
  assign cos[174]  =  12'b000111101101;     //174pi/512
  assign sin[175]  =  12'b110001111100;     //175pi/512
  assign cos[175]  =  12'b000111101000;     //175pi/512
  assign sin[176]  =  12'b110001111001;     //176pi/512
  assign cos[176]  =  12'b000111100010;     //176pi/512
  assign sin[177]  =  12'b110001110110;     //177pi/512
  assign cos[177]  =  12'b000111011101;     //177pi/512
  assign sin[178]  =  12'b110001110011;     //178pi/512
  assign cos[178]  =  12'b000111010111;     //178pi/512
  assign sin[179]  =  12'b110001110000;     //179pi/512
  assign cos[179]  =  12'b000111010010;     //179pi/512
  assign sin[180]  =  12'b110001101101;     //180pi/512
  assign cos[180]  =  12'b000111001100;     //180pi/512
  assign sin[181]  =  12'b110001101011;     //181pi/512
  assign cos[181]  =  12'b000111000110;     //181pi/512
  assign sin[182]  =  12'b110001101000;     //182pi/512
  assign cos[182]  =  12'b000111000001;     //182pi/512
  assign sin[183]  =  12'b110001100101;     //183pi/512
  assign cos[183]  =  12'b000110111011;     //183pi/512
  assign sin[184]  =  12'b110001100010;     //184pi/512
  assign cos[184]  =  12'b000110110101;     //184pi/512
  assign sin[185]  =  12'b110001100000;     //185pi/512
  assign cos[185]  =  12'b000110110000;     //185pi/512
  assign sin[186]  =  12'b110001011101;     //186pi/512
  assign cos[186]  =  12'b000110101010;     //186pi/512
  assign sin[187]  =  12'b110001011010;     //187pi/512
  assign cos[187]  =  12'b000110100100;     //187pi/512
  assign sin[188]  =  12'b110001011000;     //188pi/512
  assign cos[188]  =  12'b000110011110;     //188pi/512
  assign sin[189]  =  12'b110001010101;     //189pi/512
  assign cos[189]  =  12'b000110011001;     //189pi/512
  assign sin[190]  =  12'b110001010011;     //190pi/512
  assign cos[190]  =  12'b000110010011;     //190pi/512
  assign sin[191]  =  12'b110001010000;     //191pi/512
  assign cos[191]  =  12'b000110001101;     //191pi/512
  assign sin[192]  =  12'b110001001110;     //192pi/512
  assign cos[192]  =  12'b000110000111;     //192pi/512
  assign sin[193]  =  12'b110001001100;     //193pi/512
  assign cos[193]  =  12'b000110000010;     //193pi/512
  assign sin[194]  =  12'b110001001001;     //194pi/512
  assign cos[194]  =  12'b000101111100;     //194pi/512
  assign sin[195]  =  12'b110001000111;     //195pi/512
  assign cos[195]  =  12'b000101110110;     //195pi/512
  assign sin[196]  =  12'b110001000101;     //196pi/512
  assign cos[196]  =  12'b000101110000;     //196pi/512
  assign sin[197]  =  12'b110001000010;     //197pi/512
  assign cos[197]  =  12'b000101101010;     //197pi/512
  assign sin[198]  =  12'b110001000000;     //198pi/512
  assign cos[198]  =  12'b000101100100;     //198pi/512
  assign sin[199]  =  12'b110000111110;     //199pi/512
  assign cos[199]  =  12'b000101011110;     //199pi/512
  assign sin[200]  =  12'b110000111100;     //200pi/512
  assign cos[200]  =  12'b000101011000;     //200pi/512
  assign sin[201]  =  12'b110000111010;     //201pi/512
  assign cos[201]  =  12'b000101010011;     //201pi/512
  assign sin[202]  =  12'b110000111000;     //202pi/512
  assign cos[202]  =  12'b000101001101;     //202pi/512
  assign sin[203]  =  12'b110000110110;     //203pi/512
  assign cos[203]  =  12'b000101000111;     //203pi/512
  assign sin[204]  =  12'b110000110100;     //204pi/512
  assign cos[204]  =  12'b000101000001;     //204pi/512
  assign sin[205]  =  12'b110000110010;     //205pi/512
  assign cos[205]  =  12'b000100111011;     //205pi/512
  assign sin[206]  =  12'b110000110000;     //206pi/512
  assign cos[206]  =  12'b000100110101;     //206pi/512
  assign sin[207]  =  12'b110000101110;     //207pi/512
  assign cos[207]  =  12'b000100101111;     //207pi/512
  assign sin[208]  =  12'b110000101100;     //208pi/512
  assign cos[208]  =  12'b000100101001;     //208pi/512
  assign sin[209]  =  12'b110000101010;     //209pi/512
  assign cos[209]  =  12'b000100100011;     //209pi/512
  assign sin[210]  =  12'b110000101001;     //210pi/512
  assign cos[210]  =  12'b000100011101;     //210pi/512
  assign sin[211]  =  12'b110000100111;     //211pi/512
  assign cos[211]  =  12'b000100010111;     //211pi/512
  assign sin[212]  =  12'b110000100101;     //212pi/512
  assign cos[212]  =  12'b000100010001;     //212pi/512
  assign sin[213]  =  12'b110000100011;     //213pi/512
  assign cos[213]  =  12'b000100001011;     //213pi/512
  assign sin[214]  =  12'b110000100010;     //214pi/512
  assign cos[214]  =  12'b000100000100;     //214pi/512
  assign sin[215]  =  12'b110000100000;     //215pi/512
  assign cos[215]  =  12'b000011111110;     //215pi/512
  assign sin[216]  =  12'b110000011111;     //216pi/512
  assign cos[216]  =  12'b000011111000;     //216pi/512
  assign sin[217]  =  12'b110000011101;     //217pi/512
  assign cos[217]  =  12'b000011110010;     //217pi/512
  assign sin[218]  =  12'b110000011100;     //218pi/512
  assign cos[218]  =  12'b000011101100;     //218pi/512
  assign sin[219]  =  12'b110000011010;     //219pi/512
  assign cos[219]  =  12'b000011100110;     //219pi/512
  assign sin[220]  =  12'b110000011001;     //220pi/512
  assign cos[220]  =  12'b000011100000;     //220pi/512
  assign sin[221]  =  12'b110000011000;     //221pi/512
  assign cos[221]  =  12'b000011011010;     //221pi/512
  assign sin[222]  =  12'b110000010110;     //222pi/512
  assign cos[222]  =  12'b000011010100;     //222pi/512
  assign sin[223]  =  12'b110000010101;     //223pi/512
  assign cos[223]  =  12'b000011001101;     //223pi/512
  assign sin[224]  =  12'b110000010100;     //224pi/512
  assign cos[224]  =  12'b000011000111;     //224pi/512
  assign sin[225]  =  12'b110000010010;     //225pi/512
  assign cos[225]  =  12'b000011000001;     //225pi/512
  assign sin[226]  =  12'b110000010001;     //226pi/512
  assign cos[226]  =  12'b000010111011;     //226pi/512
  assign sin[227]  =  12'b110000010000;     //227pi/512
  assign cos[227]  =  12'b000010110101;     //227pi/512
  assign sin[228]  =  12'b110000001111;     //228pi/512
  assign cos[228]  =  12'b000010101111;     //228pi/512
  assign sin[229]  =  12'b110000001110;     //229pi/512
  assign cos[229]  =  12'b000010101000;     //229pi/512
  assign sin[230]  =  12'b110000001101;     //230pi/512
  assign cos[230]  =  12'b000010100010;     //230pi/512
  assign sin[231]  =  12'b110000001100;     //231pi/512
  assign cos[231]  =  12'b000010011100;     //231pi/512
  assign sin[232]  =  12'b110000001011;     //232pi/512
  assign cos[232]  =  12'b000010010110;     //232pi/512
  assign sin[233]  =  12'b110000001010;     //233pi/512
  assign cos[233]  =  12'b000010010000;     //233pi/512
  assign sin[234]  =  12'b110000001001;     //234pi/512
  assign cos[234]  =  12'b000010001001;     //234pi/512
  assign sin[235]  =  12'b110000001000;     //235pi/512
  assign cos[235]  =  12'b000010000011;     //235pi/512
  assign sin[236]  =  12'b110000001000;     //236pi/512
  assign cos[236]  =  12'b000001111101;     //236pi/512
  assign sin[237]  =  12'b110000000111;     //237pi/512
  assign cos[237]  =  12'b000001110111;     //237pi/512
  assign sin[238]  =  12'b110000000110;     //238pi/512
  assign cos[238]  =  12'b000001110000;     //238pi/512
  assign sin[239]  =  12'b110000000110;     //239pi/512
  assign cos[239]  =  12'b000001101010;     //239pi/512
  assign sin[240]  =  12'b110000000101;     //240pi/512
  assign cos[240]  =  12'b000001100100;     //240pi/512
  assign sin[241]  =  12'b110000000100;     //241pi/512
  assign cos[241]  =  12'b000001011110;     //241pi/512
  assign sin[242]  =  12'b110000000100;     //242pi/512
  assign cos[242]  =  12'b000001010111;     //242pi/512
  assign sin[243]  =  12'b110000000011;     //243pi/512
  assign cos[243]  =  12'b000001010001;     //243pi/512
  assign sin[244]  =  12'b110000000011;     //244pi/512
  assign cos[244]  =  12'b000001001011;     //244pi/512
  assign sin[245]  =  12'b110000000010;     //245pi/512
  assign cos[245]  =  12'b000001000101;     //245pi/512
  assign sin[246]  =  12'b110000000010;     //246pi/512
  assign cos[246]  =  12'b000000111110;     //246pi/512
  assign sin[247]  =  12'b110000000010;     //247pi/512
  assign cos[247]  =  12'b000000111000;     //247pi/512
  assign sin[248]  =  12'b110000000001;     //248pi/512
  assign cos[248]  =  12'b000000110010;     //248pi/512
  assign sin[249]  =  12'b110000000001;     //249pi/512
  assign cos[249]  =  12'b000000101011;     //249pi/512
  assign sin[250]  =  12'b110000000001;     //250pi/512
  assign cos[250]  =  12'b000000100101;     //250pi/512
  assign sin[251]  =  12'b110000000000;     //251pi/512
  assign cos[251]  =  12'b000000011111;     //251pi/512
  assign sin[252]  =  12'b110000000000;     //252pi/512
  assign cos[252]  =  12'b000000011001;     //252pi/512
  assign sin[253]  =  12'b110000000000;     //253pi/512
  assign cos[253]  =  12'b000000010010;     //253pi/512
  assign sin[254]  =  12'b110000000000;     //254pi/512
  assign cos[254]  =  12'b000000001100;     //254pi/512
  assign sin[255]  =  12'b110000000000;     //255pi/512
  assign cos[255]  =  12'b000000000110;     //255pi/512
  assign sin[256]  =  12'b110000000000;     //256pi/512
  assign cos[256]  =  12'b000000000000;     //256pi/512
  assign sin[257]  =  12'b110000000000;     //257pi/512
  assign cos[257]  =  12'b111111111010;     //257pi/512
  assign sin[258]  =  12'b110000000000;     //258pi/512
  assign cos[258]  =  12'b111111110011;     //258pi/512
  assign sin[259]  =  12'b110000000000;     //259pi/512
  assign cos[259]  =  12'b111111101101;     //259pi/512
  assign sin[260]  =  12'b110000000000;     //260pi/512
  assign cos[260]  =  12'b111111100111;     //260pi/512
  assign sin[261]  =  12'b110000000000;     //261pi/512
  assign cos[261]  =  12'b111111100001;     //261pi/512
  assign sin[262]  =  12'b110000000001;     //262pi/512
  assign cos[262]  =  12'b111111011010;     //262pi/512
  assign sin[263]  =  12'b110000000001;     //263pi/512
  assign cos[263]  =  12'b111111010100;     //263pi/512
  assign sin[264]  =  12'b110000000001;     //264pi/512
  assign cos[264]  =  12'b111111001110;     //264pi/512
  assign sin[265]  =  12'b110000000010;     //265pi/512
  assign cos[265]  =  12'b111111000111;     //265pi/512
  assign sin[266]  =  12'b110000000010;     //266pi/512
  assign cos[266]  =  12'b111111000001;     //266pi/512
  assign sin[267]  =  12'b110000000010;     //267pi/512
  assign cos[267]  =  12'b111110111011;     //267pi/512
  assign sin[268]  =  12'b110000000011;     //268pi/512
  assign cos[268]  =  12'b111110110101;     //268pi/512
  assign sin[269]  =  12'b110000000011;     //269pi/512
  assign cos[269]  =  12'b111110101110;     //269pi/512
  assign sin[270]  =  12'b110000000100;     //270pi/512
  assign cos[270]  =  12'b111110101000;     //270pi/512
  assign sin[271]  =  12'b110000000100;     //271pi/512
  assign cos[271]  =  12'b111110100010;     //271pi/512
  assign sin[272]  =  12'b110000000101;     //272pi/512
  assign cos[272]  =  12'b111110011100;     //272pi/512
  assign sin[273]  =  12'b110000000110;     //273pi/512
  assign cos[273]  =  12'b111110010101;     //273pi/512
  assign sin[274]  =  12'b110000000110;     //274pi/512
  assign cos[274]  =  12'b111110001111;     //274pi/512
  assign sin[275]  =  12'b110000000111;     //275pi/512
  assign cos[275]  =  12'b111110001001;     //275pi/512
  assign sin[276]  =  12'b110000001000;     //276pi/512
  assign cos[276]  =  12'b111110000011;     //276pi/512
  assign sin[277]  =  12'b110000001000;     //277pi/512
  assign cos[277]  =  12'b111101111100;     //277pi/512
  assign sin[278]  =  12'b110000001001;     //278pi/512
  assign cos[278]  =  12'b111101110110;     //278pi/512
  assign sin[279]  =  12'b110000001010;     //279pi/512
  assign cos[279]  =  12'b111101110000;     //279pi/512
  assign sin[280]  =  12'b110000001011;     //280pi/512
  assign cos[280]  =  12'b111101101010;     //280pi/512
  assign sin[281]  =  12'b110000001100;     //281pi/512
  assign cos[281]  =  12'b111101100100;     //281pi/512
  assign sin[282]  =  12'b110000001101;     //282pi/512
  assign cos[282]  =  12'b111101011101;     //282pi/512
  assign sin[283]  =  12'b110000001110;     //283pi/512
  assign cos[283]  =  12'b111101010111;     //283pi/512
  assign sin[284]  =  12'b110000001111;     //284pi/512
  assign cos[284]  =  12'b111101010001;     //284pi/512
  assign sin[285]  =  12'b110000010000;     //285pi/512
  assign cos[285]  =  12'b111101001011;     //285pi/512
  assign sin[286]  =  12'b110000010001;     //286pi/512
  assign cos[286]  =  12'b111101000101;     //286pi/512
  assign sin[287]  =  12'b110000010010;     //287pi/512
  assign cos[287]  =  12'b111100111110;     //287pi/512
  assign sin[288]  =  12'b110000010100;     //288pi/512
  assign cos[288]  =  12'b111100111000;     //288pi/512
  assign sin[289]  =  12'b110000010101;     //289pi/512
  assign cos[289]  =  12'b111100110010;     //289pi/512
  assign sin[290]  =  12'b110000010110;     //290pi/512
  assign cos[290]  =  12'b111100101100;     //290pi/512
  assign sin[291]  =  12'b110000011000;     //291pi/512
  assign cos[291]  =  12'b111100100110;     //291pi/512
  assign sin[292]  =  12'b110000011001;     //292pi/512
  assign cos[292]  =  12'b111100100000;     //292pi/512
  assign sin[293]  =  12'b110000011010;     //293pi/512
  assign cos[293]  =  12'b111100011010;     //293pi/512
  assign sin[294]  =  12'b110000011100;     //294pi/512
  assign cos[294]  =  12'b111100010011;     //294pi/512
  assign sin[295]  =  12'b110000011101;     //295pi/512
  assign cos[295]  =  12'b111100001101;     //295pi/512
  assign sin[296]  =  12'b110000011111;     //296pi/512
  assign cos[296]  =  12'b111100000111;     //296pi/512
  assign sin[297]  =  12'b110000100000;     //297pi/512
  assign cos[297]  =  12'b111100000001;     //297pi/512
  assign sin[298]  =  12'b110000100010;     //298pi/512
  assign cos[298]  =  12'b111011111011;     //298pi/512
  assign sin[299]  =  12'b110000100011;     //299pi/512
  assign cos[299]  =  12'b111011110101;     //299pi/512
  assign sin[300]  =  12'b110000100101;     //300pi/512
  assign cos[300]  =  12'b111011101111;     //300pi/512
  assign sin[301]  =  12'b110000100111;     //301pi/512
  assign cos[301]  =  12'b111011101001;     //301pi/512
  assign sin[302]  =  12'b110000101001;     //302pi/512
  assign cos[302]  =  12'b111011100011;     //302pi/512
  assign sin[303]  =  12'b110000101010;     //303pi/512
  assign cos[303]  =  12'b111011011101;     //303pi/512
  assign sin[304]  =  12'b110000101100;     //304pi/512
  assign cos[304]  =  12'b111011010111;     //304pi/512
  assign sin[305]  =  12'b110000101110;     //305pi/512
  assign cos[305]  =  12'b111011010001;     //305pi/512
  assign sin[306]  =  12'b110000110000;     //306pi/512
  assign cos[306]  =  12'b111011001011;     //306pi/512
  assign sin[307]  =  12'b110000110010;     //307pi/512
  assign cos[307]  =  12'b111011000101;     //307pi/512
  assign sin[308]  =  12'b110000110100;     //308pi/512
  assign cos[308]  =  12'b111010111111;     //308pi/512
  assign sin[309]  =  12'b110000110110;     //309pi/512
  assign cos[309]  =  12'b111010111001;     //309pi/512
  assign sin[310]  =  12'b110000111000;     //310pi/512
  assign cos[310]  =  12'b111010110011;     //310pi/512
  assign sin[311]  =  12'b110000111010;     //311pi/512
  assign cos[311]  =  12'b111010101101;     //311pi/512
  assign sin[312]  =  12'b110000111100;     //312pi/512
  assign cos[312]  =  12'b111010100111;     //312pi/512
  assign sin[313]  =  12'b110000111110;     //313pi/512
  assign cos[313]  =  12'b111010100001;     //313pi/512
  assign sin[314]  =  12'b110001000000;     //314pi/512
  assign cos[314]  =  12'b111010011011;     //314pi/512
  assign sin[315]  =  12'b110001000010;     //315pi/512
  assign cos[315]  =  12'b111010010101;     //315pi/512
  assign sin[316]  =  12'b110001000101;     //316pi/512
  assign cos[316]  =  12'b111010001111;     //316pi/512
  assign sin[317]  =  12'b110001000111;     //317pi/512
  assign cos[317]  =  12'b111010001010;     //317pi/512
  assign sin[318]  =  12'b110001001001;     //318pi/512
  assign cos[318]  =  12'b111010000100;     //318pi/512
  assign sin[319]  =  12'b110001001100;     //319pi/512
  assign cos[319]  =  12'b111001111110;     //319pi/512
  assign sin[320]  =  12'b110001001110;     //320pi/512
  assign cos[320]  =  12'b111001111000;     //320pi/512
  assign sin[321]  =  12'b110001010000;     //321pi/512
  assign cos[321]  =  12'b111001110010;     //321pi/512
  assign sin[322]  =  12'b110001010011;     //322pi/512
  assign cos[322]  =  12'b111001101101;     //322pi/512
  assign sin[323]  =  12'b110001010101;     //323pi/512
  assign cos[323]  =  12'b111001100111;     //323pi/512
  assign sin[324]  =  12'b110001011000;     //324pi/512
  assign cos[324]  =  12'b111001100001;     //324pi/512
  assign sin[325]  =  12'b110001011010;     //325pi/512
  assign cos[325]  =  12'b111001011011;     //325pi/512
  assign sin[326]  =  12'b110001011101;     //326pi/512
  assign cos[326]  =  12'b111001010110;     //326pi/512
  assign sin[327]  =  12'b110001100000;     //327pi/512
  assign cos[327]  =  12'b111001010000;     //327pi/512
  assign sin[328]  =  12'b110001100010;     //328pi/512
  assign cos[328]  =  12'b111001001010;     //328pi/512
  assign sin[329]  =  12'b110001100101;     //329pi/512
  assign cos[329]  =  12'b111001000101;     //329pi/512
  assign sin[330]  =  12'b110001101000;     //330pi/512
  assign cos[330]  =  12'b111000111111;     //330pi/512
  assign sin[331]  =  12'b110001101011;     //331pi/512
  assign cos[331]  =  12'b111000111001;     //331pi/512
  assign sin[332]  =  12'b110001101101;     //332pi/512
  assign cos[332]  =  12'b111000110100;     //332pi/512
  assign sin[333]  =  12'b110001110000;     //333pi/512
  assign cos[333]  =  12'b111000101110;     //333pi/512
  assign sin[334]  =  12'b110001110011;     //334pi/512
  assign cos[334]  =  12'b111000101000;     //334pi/512
  assign sin[335]  =  12'b110001110110;     //335pi/512
  assign cos[335]  =  12'b111000100011;     //335pi/512
  assign sin[336]  =  12'b110001111001;     //336pi/512
  assign cos[336]  =  12'b111000011101;     //336pi/512
  assign sin[337]  =  12'b110001111100;     //337pi/512
  assign cos[337]  =  12'b111000011000;     //337pi/512
  assign sin[338]  =  12'b110001111111;     //338pi/512
  assign cos[338]  =  12'b111000010010;     //338pi/512
  assign sin[339]  =  12'b110010000010;     //339pi/512
  assign cos[339]  =  12'b111000001101;     //339pi/512
  assign sin[340]  =  12'b110010000101;     //340pi/512
  assign cos[340]  =  12'b111000000111;     //340pi/512
  assign sin[341]  =  12'b110010001000;     //341pi/512
  assign cos[341]  =  12'b111000000010;     //341pi/512
  assign sin[342]  =  12'b110010001011;     //342pi/512
  assign cos[342]  =  12'b110111111100;     //342pi/512
  assign sin[343]  =  12'b110010001110;     //343pi/512
  assign cos[343]  =  12'b110111110111;     //343pi/512
  assign sin[344]  =  12'b110010010010;     //344pi/512
  assign cos[344]  =  12'b110111110010;     //344pi/512
  assign sin[345]  =  12'b110010010101;     //345pi/512
  assign cos[345]  =  12'b110111101100;     //345pi/512
  assign sin[346]  =  12'b110010011000;     //346pi/512
  assign cos[346]  =  12'b110111100111;     //346pi/512
  assign sin[347]  =  12'b110010011100;     //347pi/512
  assign cos[347]  =  12'b110111100001;     //347pi/512
  assign sin[348]  =  12'b110010011111;     //348pi/512
  assign cos[348]  =  12'b110111011100;     //348pi/512
  assign sin[349]  =  12'b110010100010;     //349pi/512
  assign cos[349]  =  12'b110111010111;     //349pi/512
  assign sin[350]  =  12'b110010100110;     //350pi/512
  assign cos[350]  =  12'b110111010010;     //350pi/512
  assign sin[351]  =  12'b110010101001;     //351pi/512
  assign cos[351]  =  12'b110111001100;     //351pi/512
  assign sin[352]  =  12'b110010101101;     //352pi/512
  assign cos[352]  =  12'b110111000111;     //352pi/512
  assign sin[353]  =  12'b110010110000;     //353pi/512
  assign cos[353]  =  12'b110111000010;     //353pi/512
  assign sin[354]  =  12'b110010110100;     //354pi/512
  assign cos[354]  =  12'b110110111101;     //354pi/512
  assign sin[355]  =  12'b110010110111;     //355pi/512
  assign cos[355]  =  12'b110110111000;     //355pi/512
  assign sin[356]  =  12'b110010111011;     //356pi/512
  assign cos[356]  =  12'b110110110010;     //356pi/512
  assign sin[357]  =  12'b110010111110;     //357pi/512
  assign cos[357]  =  12'b110110101101;     //357pi/512
  assign sin[358]  =  12'b110011000010;     //358pi/512
  assign cos[358]  =  12'b110110101000;     //358pi/512
  assign sin[359]  =  12'b110011000110;     //359pi/512
  assign cos[359]  =  12'b110110100011;     //359pi/512
  assign sin[360]  =  12'b110011001010;     //360pi/512
  assign cos[360]  =  12'b110110011110;     //360pi/512
  assign sin[361]  =  12'b110011001101;     //361pi/512
  assign cos[361]  =  12'b110110011001;     //361pi/512
  assign sin[362]  =  12'b110011010001;     //362pi/512
  assign cos[362]  =  12'b110110010100;     //362pi/512
  assign sin[363]  =  12'b110011010101;     //363pi/512
  assign cos[363]  =  12'b110110001111;     //363pi/512
  assign sin[364]  =  12'b110011011001;     //364pi/512
  assign cos[364]  =  12'b110110001010;     //364pi/512
  assign sin[365]  =  12'b110011011101;     //365pi/512
  assign cos[365]  =  12'b110110000101;     //365pi/512
  assign sin[366]  =  12'b110011100001;     //366pi/512
  assign cos[366]  =  12'b110110000000;     //366pi/512
  assign sin[367]  =  12'b110011100100;     //367pi/512
  assign cos[367]  =  12'b110101111011;     //367pi/512
  assign sin[368]  =  12'b110011101000;     //368pi/512
  assign cos[368]  =  12'b110101110110;     //368pi/512
  assign sin[369]  =  12'b110011101100;     //369pi/512
  assign cos[369]  =  12'b110101110010;     //369pi/512
  assign sin[370]  =  12'b110011110000;     //370pi/512
  assign cos[370]  =  12'b110101101101;     //370pi/512
  assign sin[371]  =  12'b110011110101;     //371pi/512
  assign cos[371]  =  12'b110101101000;     //371pi/512
  assign sin[372]  =  12'b110011111001;     //372pi/512
  assign cos[372]  =  12'b110101100011;     //372pi/512
  assign sin[373]  =  12'b110011111101;     //373pi/512
  assign cos[373]  =  12'b110101011110;     //373pi/512
  assign sin[374]  =  12'b110100000001;     //374pi/512
  assign cos[374]  =  12'b110101011010;     //374pi/512
  assign sin[375]  =  12'b110100000101;     //375pi/512
  assign cos[375]  =  12'b110101010101;     //375pi/512
  assign sin[376]  =  12'b110100001001;     //376pi/512
  assign cos[376]  =  12'b110101010000;     //376pi/512
  assign sin[377]  =  12'b110100001101;     //377pi/512
  assign cos[377]  =  12'b110101001100;     //377pi/512
  assign sin[378]  =  12'b110100010010;     //378pi/512
  assign cos[378]  =  12'b110101000111;     //378pi/512
  assign sin[379]  =  12'b110100010110;     //379pi/512
  assign cos[379]  =  12'b110101000010;     //379pi/512
  assign sin[380]  =  12'b110100011010;     //380pi/512
  assign cos[380]  =  12'b110100111110;     //380pi/512
  assign sin[381]  =  12'b110100011111;     //381pi/512
  assign cos[381]  =  12'b110100111001;     //381pi/512
  assign sin[382]  =  12'b110100100011;     //382pi/512
  assign cos[382]  =  12'b110100110101;     //382pi/512
  assign sin[383]  =  12'b110100100111;     //383pi/512
  assign cos[383]  =  12'b110100110000;     //383pi/512
  assign sin[384]  =  12'b110100101100;     //384pi/512
  assign cos[384]  =  12'b110100101100;     //384pi/512
  assign sin[385]  =  12'b110100110000;     //385pi/512
  assign cos[385]  =  12'b110100100111;     //385pi/512
  assign sin[386]  =  12'b110100110101;     //386pi/512
  assign cos[386]  =  12'b110100100011;     //386pi/512
  assign sin[387]  =  12'b110100111001;     //387pi/512
  assign cos[387]  =  12'b110100011111;     //387pi/512
  assign sin[388]  =  12'b110100111110;     //388pi/512
  assign cos[388]  =  12'b110100011010;     //388pi/512
  assign sin[389]  =  12'b110101000010;     //389pi/512
  assign cos[389]  =  12'b110100010110;     //389pi/512
  assign sin[390]  =  12'b110101000111;     //390pi/512
  assign cos[390]  =  12'b110100010010;     //390pi/512
  assign sin[391]  =  12'b110101001100;     //391pi/512
  assign cos[391]  =  12'b110100001101;     //391pi/512
  assign sin[392]  =  12'b110101010000;     //392pi/512
  assign cos[392]  =  12'b110100001001;     //392pi/512
  assign sin[393]  =  12'b110101010101;     //393pi/512
  assign cos[393]  =  12'b110100000101;     //393pi/512
  assign sin[394]  =  12'b110101011010;     //394pi/512
  assign cos[394]  =  12'b110100000001;     //394pi/512
  assign sin[395]  =  12'b110101011110;     //395pi/512
  assign cos[395]  =  12'b110011111101;     //395pi/512
  assign sin[396]  =  12'b110101100011;     //396pi/512
  assign cos[396]  =  12'b110011111001;     //396pi/512
  assign sin[397]  =  12'b110101101000;     //397pi/512
  assign cos[397]  =  12'b110011110101;     //397pi/512
  assign sin[398]  =  12'b110101101101;     //398pi/512
  assign cos[398]  =  12'b110011110000;     //398pi/512
  assign sin[399]  =  12'b110101110010;     //399pi/512
  assign cos[399]  =  12'b110011101100;     //399pi/512
  assign sin[400]  =  12'b110101110110;     //400pi/512
  assign cos[400]  =  12'b110011101000;     //400pi/512
  assign sin[401]  =  12'b110101111011;     //401pi/512
  assign cos[401]  =  12'b110011100100;     //401pi/512
  assign sin[402]  =  12'b110110000000;     //402pi/512
  assign cos[402]  =  12'b110011100001;     //402pi/512
  assign sin[403]  =  12'b110110000101;     //403pi/512
  assign cos[403]  =  12'b110011011101;     //403pi/512
  assign sin[404]  =  12'b110110001010;     //404pi/512
  assign cos[404]  =  12'b110011011001;     //404pi/512
  assign sin[405]  =  12'b110110001111;     //405pi/512
  assign cos[405]  =  12'b110011010101;     //405pi/512
  assign sin[406]  =  12'b110110010100;     //406pi/512
  assign cos[406]  =  12'b110011010001;     //406pi/512
  assign sin[407]  =  12'b110110011001;     //407pi/512
  assign cos[407]  =  12'b110011001101;     //407pi/512
  assign sin[408]  =  12'b110110011110;     //408pi/512
  assign cos[408]  =  12'b110011001010;     //408pi/512
  assign sin[409]  =  12'b110110100011;     //409pi/512
  assign cos[409]  =  12'b110011000110;     //409pi/512
  assign sin[410]  =  12'b110110101000;     //410pi/512
  assign cos[410]  =  12'b110011000010;     //410pi/512
  assign sin[411]  =  12'b110110101101;     //411pi/512
  assign cos[411]  =  12'b110010111110;     //411pi/512
  assign sin[412]  =  12'b110110110010;     //412pi/512
  assign cos[412]  =  12'b110010111011;     //412pi/512
  assign sin[413]  =  12'b110110111000;     //413pi/512
  assign cos[413]  =  12'b110010110111;     //413pi/512
  assign sin[414]  =  12'b110110111101;     //414pi/512
  assign cos[414]  =  12'b110010110100;     //414pi/512
  assign sin[415]  =  12'b110111000010;     //415pi/512
  assign cos[415]  =  12'b110010110000;     //415pi/512
  assign sin[416]  =  12'b110111000111;     //416pi/512
  assign cos[416]  =  12'b110010101101;     //416pi/512
  assign sin[417]  =  12'b110111001100;     //417pi/512
  assign cos[417]  =  12'b110010101001;     //417pi/512
  assign sin[418]  =  12'b110111010010;     //418pi/512
  assign cos[418]  =  12'b110010100110;     //418pi/512
  assign sin[419]  =  12'b110111010111;     //419pi/512
  assign cos[419]  =  12'b110010100010;     //419pi/512
  assign sin[420]  =  12'b110111011100;     //420pi/512
  assign cos[420]  =  12'b110010011111;     //420pi/512
  assign sin[421]  =  12'b110111100001;     //421pi/512
  assign cos[421]  =  12'b110010011100;     //421pi/512
  assign sin[422]  =  12'b110111100111;     //422pi/512
  assign cos[422]  =  12'b110010011000;     //422pi/512
  assign sin[423]  =  12'b110111101100;     //423pi/512
  assign cos[423]  =  12'b110010010101;     //423pi/512
  assign sin[424]  =  12'b110111110010;     //424pi/512
  assign cos[424]  =  12'b110010010010;     //424pi/512
  assign sin[425]  =  12'b110111110111;     //425pi/512
  assign cos[425]  =  12'b110010001110;     //425pi/512
  assign sin[426]  =  12'b110111111100;     //426pi/512
  assign cos[426]  =  12'b110010001011;     //426pi/512
  assign sin[427]  =  12'b111000000010;     //427pi/512
  assign cos[427]  =  12'b110010001000;     //427pi/512
  assign sin[428]  =  12'b111000000111;     //428pi/512
  assign cos[428]  =  12'b110010000101;     //428pi/512
  assign sin[429]  =  12'b111000001101;     //429pi/512
  assign cos[429]  =  12'b110010000010;     //429pi/512
  assign sin[430]  =  12'b111000010010;     //430pi/512
  assign cos[430]  =  12'b110001111111;     //430pi/512
  assign sin[431]  =  12'b111000011000;     //431pi/512
  assign cos[431]  =  12'b110001111100;     //431pi/512
  assign sin[432]  =  12'b111000011101;     //432pi/512
  assign cos[432]  =  12'b110001111001;     //432pi/512
  assign sin[433]  =  12'b111000100011;     //433pi/512
  assign cos[433]  =  12'b110001110110;     //433pi/512
  assign sin[434]  =  12'b111000101000;     //434pi/512
  assign cos[434]  =  12'b110001110011;     //434pi/512
  assign sin[435]  =  12'b111000101110;     //435pi/512
  assign cos[435]  =  12'b110001110000;     //435pi/512
  assign sin[436]  =  12'b111000110100;     //436pi/512
  assign cos[436]  =  12'b110001101101;     //436pi/512
  assign sin[437]  =  12'b111000111001;     //437pi/512
  assign cos[437]  =  12'b110001101011;     //437pi/512
  assign sin[438]  =  12'b111000111111;     //438pi/512
  assign cos[438]  =  12'b110001101000;     //438pi/512
  assign sin[439]  =  12'b111001000101;     //439pi/512
  assign cos[439]  =  12'b110001100101;     //439pi/512
  assign sin[440]  =  12'b111001001010;     //440pi/512
  assign cos[440]  =  12'b110001100010;     //440pi/512
  assign sin[441]  =  12'b111001010000;     //441pi/512
  assign cos[441]  =  12'b110001100000;     //441pi/512
  assign sin[442]  =  12'b111001010110;     //442pi/512
  assign cos[442]  =  12'b110001011101;     //442pi/512
  assign sin[443]  =  12'b111001011011;     //443pi/512
  assign cos[443]  =  12'b110001011010;     //443pi/512
  assign sin[444]  =  12'b111001100001;     //444pi/512
  assign cos[444]  =  12'b110001011000;     //444pi/512
  assign sin[445]  =  12'b111001100111;     //445pi/512
  assign cos[445]  =  12'b110001010101;     //445pi/512
  assign sin[446]  =  12'b111001101101;     //446pi/512
  assign cos[446]  =  12'b110001010011;     //446pi/512
  assign sin[447]  =  12'b111001110010;     //447pi/512
  assign cos[447]  =  12'b110001010000;     //447pi/512
  assign sin[448]  =  12'b111001111000;     //448pi/512
  assign cos[448]  =  12'b110001001110;     //448pi/512
  assign sin[449]  =  12'b111001111110;     //449pi/512
  assign cos[449]  =  12'b110001001100;     //449pi/512
  assign sin[450]  =  12'b111010000100;     //450pi/512
  assign cos[450]  =  12'b110001001001;     //450pi/512
  assign sin[451]  =  12'b111010001010;     //451pi/512
  assign cos[451]  =  12'b110001000111;     //451pi/512
  assign sin[452]  =  12'b111010001111;     //452pi/512
  assign cos[452]  =  12'b110001000101;     //452pi/512
  assign sin[453]  =  12'b111010010101;     //453pi/512
  assign cos[453]  =  12'b110001000010;     //453pi/512
  assign sin[454]  =  12'b111010011011;     //454pi/512
  assign cos[454]  =  12'b110001000000;     //454pi/512
  assign sin[455]  =  12'b111010100001;     //455pi/512
  assign cos[455]  =  12'b110000111110;     //455pi/512
  assign sin[456]  =  12'b111010100111;     //456pi/512
  assign cos[456]  =  12'b110000111100;     //456pi/512
  assign sin[457]  =  12'b111010101101;     //457pi/512
  assign cos[457]  =  12'b110000111010;     //457pi/512
  assign sin[458]  =  12'b111010110011;     //458pi/512
  assign cos[458]  =  12'b110000111000;     //458pi/512
  assign sin[459]  =  12'b111010111001;     //459pi/512
  assign cos[459]  =  12'b110000110110;     //459pi/512
  assign sin[460]  =  12'b111010111111;     //460pi/512
  assign cos[460]  =  12'b110000110100;     //460pi/512
  assign sin[461]  =  12'b111011000101;     //461pi/512
  assign cos[461]  =  12'b110000110010;     //461pi/512
  assign sin[462]  =  12'b111011001011;     //462pi/512
  assign cos[462]  =  12'b110000110000;     //462pi/512
  assign sin[463]  =  12'b111011010001;     //463pi/512
  assign cos[463]  =  12'b110000101110;     //463pi/512
  assign sin[464]  =  12'b111011010111;     //464pi/512
  assign cos[464]  =  12'b110000101100;     //464pi/512
  assign sin[465]  =  12'b111011011101;     //465pi/512
  assign cos[465]  =  12'b110000101010;     //465pi/512
  assign sin[466]  =  12'b111011100011;     //466pi/512
  assign cos[466]  =  12'b110000101001;     //466pi/512
  assign sin[467]  =  12'b111011101001;     //467pi/512
  assign cos[467]  =  12'b110000100111;     //467pi/512
  assign sin[468]  =  12'b111011101111;     //468pi/512
  assign cos[468]  =  12'b110000100101;     //468pi/512
  assign sin[469]  =  12'b111011110101;     //469pi/512
  assign cos[469]  =  12'b110000100011;     //469pi/512
  assign sin[470]  =  12'b111011111011;     //470pi/512
  assign cos[470]  =  12'b110000100010;     //470pi/512
  assign sin[471]  =  12'b111100000001;     //471pi/512
  assign cos[471]  =  12'b110000100000;     //471pi/512
  assign sin[472]  =  12'b111100000111;     //472pi/512
  assign cos[472]  =  12'b110000011111;     //472pi/512
  assign sin[473]  =  12'b111100001101;     //473pi/512
  assign cos[473]  =  12'b110000011101;     //473pi/512
  assign sin[474]  =  12'b111100010011;     //474pi/512
  assign cos[474]  =  12'b110000011100;     //474pi/512
  assign sin[475]  =  12'b111100011010;     //475pi/512
  assign cos[475]  =  12'b110000011010;     //475pi/512
  assign sin[476]  =  12'b111100100000;     //476pi/512
  assign cos[476]  =  12'b110000011001;     //476pi/512
  assign sin[477]  =  12'b111100100110;     //477pi/512
  assign cos[477]  =  12'b110000011000;     //477pi/512
  assign sin[478]  =  12'b111100101100;     //478pi/512
  assign cos[478]  =  12'b110000010110;     //478pi/512
  assign sin[479]  =  12'b111100110010;     //479pi/512
  assign cos[479]  =  12'b110000010101;     //479pi/512
  assign sin[480]  =  12'b111100111000;     //480pi/512
  assign cos[480]  =  12'b110000010100;     //480pi/512
  assign sin[481]  =  12'b111100111110;     //481pi/512
  assign cos[481]  =  12'b110000010010;     //481pi/512
  assign sin[482]  =  12'b111101000101;     //482pi/512
  assign cos[482]  =  12'b110000010001;     //482pi/512
  assign sin[483]  =  12'b111101001011;     //483pi/512
  assign cos[483]  =  12'b110000010000;     //483pi/512
  assign sin[484]  =  12'b111101010001;     //484pi/512
  assign cos[484]  =  12'b110000001111;     //484pi/512
  assign sin[485]  =  12'b111101010111;     //485pi/512
  assign cos[485]  =  12'b110000001110;     //485pi/512
  assign sin[486]  =  12'b111101011101;     //486pi/512
  assign cos[486]  =  12'b110000001101;     //486pi/512
  assign sin[487]  =  12'b111101100100;     //487pi/512
  assign cos[487]  =  12'b110000001100;     //487pi/512
  assign sin[488]  =  12'b111101101010;     //488pi/512
  assign cos[488]  =  12'b110000001011;     //488pi/512
  assign sin[489]  =  12'b111101110000;     //489pi/512
  assign cos[489]  =  12'b110000001010;     //489pi/512
  assign sin[490]  =  12'b111101110110;     //490pi/512
  assign cos[490]  =  12'b110000001001;     //490pi/512
  assign sin[491]  =  12'b111101111100;     //491pi/512
  assign cos[491]  =  12'b110000001000;     //491pi/512
  assign sin[492]  =  12'b111110000011;     //492pi/512
  assign cos[492]  =  12'b110000001000;     //492pi/512
  assign sin[493]  =  12'b111110001001;     //493pi/512
  assign cos[493]  =  12'b110000000111;     //493pi/512
  assign sin[494]  =  12'b111110001111;     //494pi/512
  assign cos[494]  =  12'b110000000110;     //494pi/512
  assign sin[495]  =  12'b111110010101;     //495pi/512
  assign cos[495]  =  12'b110000000110;     //495pi/512
  assign sin[496]  =  12'b111110011100;     //496pi/512
  assign cos[496]  =  12'b110000000101;     //496pi/512
  assign sin[497]  =  12'b111110100010;     //497pi/512
  assign cos[497]  =  12'b110000000100;     //497pi/512
  assign sin[498]  =  12'b111110101000;     //498pi/512
  assign cos[498]  =  12'b110000000100;     //498pi/512
  assign sin[499]  =  12'b111110101110;     //499pi/512
  assign cos[499]  =  12'b110000000011;     //499pi/512
  assign sin[500]  =  12'b111110110101;     //500pi/512
  assign cos[500]  =  12'b110000000011;     //500pi/512
  assign sin[501]  =  12'b111110111011;     //501pi/512
  assign cos[501]  =  12'b110000000010;     //501pi/512
  assign sin[502]  =  12'b111111000001;     //502pi/512
  assign cos[502]  =  12'b110000000010;     //502pi/512
  assign sin[503]  =  12'b111111000111;     //503pi/512
  assign cos[503]  =  12'b110000000010;     //503pi/512
  assign sin[504]  =  12'b111111001110;     //504pi/512
  assign cos[504]  =  12'b110000000001;     //504pi/512
  assign sin[505]  =  12'b111111010100;     //505pi/512
  assign cos[505]  =  12'b110000000001;     //505pi/512
  assign sin[506]  =  12'b111111011010;     //506pi/512
  assign cos[506]  =  12'b110000000001;     //506pi/512
  assign sin[507]  =  12'b111111100001;     //507pi/512
  assign cos[507]  =  12'b110000000000;     //507pi/512
  assign sin[508]  =  12'b111111100111;     //508pi/512
  assign cos[508]  =  12'b110000000000;     //508pi/512
  assign sin[509]  =  12'b111111101101;     //509pi/512
  assign cos[509]  =  12'b110000000000;     //509pi/512
  assign sin[510]  =  12'b111111110011;     //510pi/512
  assign cos[510]  =  12'b110000000000;     //510pi/512
  assign sin[511]  =  12'b111111111010;     //511pi/512
  assign cos[511]  =  12'b110000000000;     //511pi/512

endmodule