module  RAM #(parameter bit_width=29, N = 16, SIZE = 4)(
    input                              clk,rst_n,
    
    input                              load_data,
    input              [SIZE:       0] invert_adr,
    input       signed [bit_width-1:0] Re_i1,
    input       signed [bit_width-1:0] Im_i1,

    input                               en_wr,
    input              [SIZE:       0]  wr_ptr,
    input       signed [bit_width-1:0]  Re_i2,
    input       signed [bit_width-1:0]  Im_i2,

    
    input              [SIZE:       0]  rd_ptr,
    input                               en_rd, 
    input                               finish_FFT,
    input                               done_all, 
    input              [10          :0] rd_angle_ptr,
    
    output reg  signed [bit_width-1:0]  Re_o1,
    output reg  signed [bit_width-1:0]  Im_o1,
    output reg  signed [bit_width-1:0]  Re_o2,
    output reg  signed [bit_width-1:0]  Im_o2,
    output reg                          en_add,       

    output reg  signed [bit_width-1:0]  Re_o,
    output reg  signed [bit_width-1:0]  Im_o,

    output  reg signed [13         :0]  cos_data,
    output  reg signed [13         :0]  sin_data,
    
    output reg                          en_o
 );

    reg  signed [bit_width-1:0]   x_real_i;
    reg  signed [bit_width-1:0]   y_real_i;
    reg         [SIZE:       0]   index_wr ;


    reg  signed  [bit_width-1:0]  mem_Re  [N-1:0];
    reg  signed  [bit_width-1:0]  mem_Im  [N-1:0];

    reg  signed  [bit_width-1:0]  Re_o_temp;
    reg  signed  [bit_width-1:0]  Im_o_temp;

    reg  signed  [bit_width-1:0]  Re_o1_temp;
    reg  signed  [bit_width-1:0]  Im_o1_temp;
    
    reg                           en_o_temp;
    
    reg  en_o_1, en_o_2;
    reg  en_wr_mem;
    
    reg [1:0] state;
    reg [1:0] state2;

    reg signed [13:0]  cos  [255:0];
    reg signed [13:0]  sin  [255:0];

  //  assign en_add = en_o_2;

    localparam 
          FIRST_OUT = 2'b01,
          SEC_OUT   = 2'b10;
    localparam
          PROCESS   = 2'b01,
          FINISH    = 2'b10;  
    //--------------------handle choose out put------------------------------  
        always @(posedge clk or negedge rst_n) begin
            if (!rst_n) begin
                state          <= FIRST_OUT;
                en_o_1         <= 1'b0;  
                en_o_2         <= 1'b0;
            end else begin
                case (state)
                  FIRST_OUT  : begin
                    if (en_rd) begin
                        en_o_1         <= 1'b1;  
                        en_o_2         <= 1'b0;
                        state          <= SEC_OUT;
                    end 
                    end
                  SEC_OUT: begin
                        en_o_2         <= 1'b1;
                        en_o_1         <= 1'b0;
                        state     <= FIRST_OUT;
                  end
                    default: state     <= FIRST_OUT;
                endcase
            end
        end
        always @(posedge clk) begin
                if (en_o_1) begin
                Re_o1_temp       <= Re_o_temp;
                Im_o1_temp       <= Im_o_temp;
                end
        end 
       always @(*) begin
                if (en_o_2) begin
                    Re_o2  <= Re_o_temp;
                    Im_o2  <= Im_o_temp;
                    Re_o1  <= Re_o1_temp;
                    Im_o1  <= Im_o1_temp;
                    en_add <= 1'b1;
                end else en_add <= 1'b0;
        end  
    //--------------------handle out put------------------------------  
        always @(posedge clk or negedge rst_n) begin
            if (!rst_n) begin
                state2   <=   PROCESS;
                en_o    <= 0; 
            end else begin
                case (state2)
                  PROCESS  : begin
                    if (finish_FFT) state2   <= FINISH;   
                    en_o    <= 0;   
                    end
                  FINISH: begin
                        Re_o      <= Re_o_temp;
                        Im_o      <= Im_o_temp;
                        en_o      <= en_o_temp;
                    if (done_all) 
                        state2     <= PROCESS;
                  end
                    default: state2     <= PROCESS;
                endcase
            end
        end
    //------------------------handle read write from MEM----------------------------
        always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            Re_o_temp      <= 0;
            Im_o_temp      <= 0;
            en_o_temp      <= 0;
        end else begin
             if (en_rd) begin
                  Re_o_temp             <= mem_Re[rd_ptr];
                  Im_o_temp             <= mem_Im[rd_ptr];
                  en_o_temp             <= 1'b1;
             end else  en_o_temp        <= 0;
             if (en_wr_mem) begin
                  mem_Re[index_wr] <= x_real_i;
                  mem_Im[index_wr] <= y_real_i;    
            end
        end
        end
    //------------------------handle load initial data to MEM--------------------------
        always @(posedge clk or negedge rst_n) begin
            if (!rst_n) begin
                en_wr_mem <= 1'b0;
            end else if (load_data) begin
                x_real_i  <= Re_i1;
                y_real_i  <= Im_i1;
                index_wr  <= invert_adr; 
                en_wr_mem <= 1'b1;
            end else if (en_wr) begin
                x_real_i  <= Re_i2;
                y_real_i  <= Im_i2;
                index_wr  <= wr_ptr; 
                en_wr_mem <= 1'b1;
            end else en_wr_mem <= 1'b0;
        end

    //--------------------------------handle reaf tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd ) begin
                  cos_data         <= cos   [rd_angle_ptr];
                  sin_data         <= sin   [rd_angle_ptr];
             end
        end

//------------------------ROM-------------------------------------------------------
initial begin
   sin[0]  =  14'b00000000000000;     //0pi/128
   cos[0]  =  14'b01000000000000;     //0pi/128
   sin[1]  =  14'b11111110011011;     //1pi/128
   cos[1]  =  14'b00111111111110;     //1pi/128
   sin[2]  =  14'b11111100110111;     //2pi/128
   cos[2]  =  14'b00111111111011;     //2pi/128
   sin[3]  =  14'b11111011010011;     //3pi/128
   cos[3]  =  14'b00111111110100;     //3pi/128
   sin[4]  =  14'b11111001101111;     //4pi/128
   cos[4]  =  14'b00111111101100;     //4pi/128
   sin[5]  =  14'b11111000001011;     //5pi/128
   cos[5]  =  14'b00111111100001;     //5pi/128
   sin[6]  =  14'b11110110100111;     //6pi/128
   cos[6]  =  14'b00111111010011;     //6pi/128
   sin[7]  =  14'b11110101000100;     //7pi/128
   cos[7]  =  14'b00111111000011;     //7pi/128
   sin[8]  =  14'b11110011100001;     //8pi/128
   cos[8]  =  14'b00111110110001;     //8pi/128
   sin[9]  =  14'b11110001111111;     //9pi/128
   cos[9]  =  14'b00111110011100;     //9pi/128
   sin[10]  =  14'b11110000011101;     //10pi/128
   cos[10]  =  14'b00111110000101;     //10pi/128
   sin[11]  =  14'b11101110111100;     //11pi/128
   cos[11]  =  14'b00111101101011;     //11pi/128
   sin[12]  =  14'b11101101011011;     //12pi/128
   cos[12]  =  14'b00111101001111;     //12pi/128
   sin[13]  =  14'b11101011111011;     //13pi/128
   cos[13]  =  14'b00111100110001;     //13pi/128
   sin[14]  =  14'b11101010011100;     //14pi/128
   cos[14]  =  14'b00111100010000;     //14pi/128
   sin[15]  =  14'b11101000111110;     //15pi/128
   cos[15]  =  14'b00111011101101;     //15pi/128
   sin[16]  =  14'b11100111100001;     //16pi/128
   cos[16]  =  14'b00111011001000;     //16pi/128
   sin[17]  =  14'b11100110000100;     //17pi/128
   cos[17]  =  14'b00111010100000;     //17pi/128
   sin[18]  =  14'b11100100101001;     //18pi/128
   cos[18]  =  14'b00111001110110;     //18pi/128
   sin[19]  =  14'b11100011001110;     //19pi/128
   cos[19]  =  14'b00111001001010;     //19pi/128
   sin[20]  =  14'b11100001110101;     //20pi/128
   cos[20]  =  14'b00111000011100;     //20pi/128
   sin[21]  =  14'b11100000011101;     //21pi/128
   cos[21]  =  14'b00110111101011;     //21pi/128
   sin[22]  =  14'b11011111000110;     //22pi/128
   cos[22]  =  14'b00110110111001;     //22pi/128
   sin[23]  =  14'b11011101110001;     //23pi/128
   cos[23]  =  14'b00110110000100;     //23pi/128
   sin[24]  =  14'b11011100011100;     //24pi/128
   cos[24]  =  14'b00110101001101;     //24pi/128
   sin[25]  =  14'b11011011001001;     //25pi/128
   cos[25]  =  14'b00110100010100;     //25pi/128
   sin[26]  =  14'b11011001111000;     //26pi/128
   cos[26]  =  14'b00110011011001;     //26pi/128
   sin[27]  =  14'b11011000101000;     //27pi/128
   cos[27]  =  14'b00110010011101;     //27pi/128
   sin[28]  =  14'b11010111011010;     //28pi/128
   cos[28]  =  14'b00110001011110;     //28pi/128
   sin[29]  =  14'b11010110001101;     //29pi/128
   cos[29]  =  14'b00110000011101;     //29pi/128
   sin[30]  =  14'b11010101000001;     //30pi/128
   cos[30]  =  14'b00101111011010;     //30pi/128
   sin[31]  =  14'b11010011111000;     //31pi/128
   cos[31]  =  14'b00101110010110;     //31pi/128
   sin[32]  =  14'b11010010110000;     //32pi/128
   cos[32]  =  14'b00101101010000;     //32pi/128
   sin[33]  =  14'b11010001101001;     //33pi/128
   cos[33]  =  14'b00101100001000;     //33pi/128
   sin[34]  =  14'b11010000100101;     //34pi/128
   cos[34]  =  14'b00101010111110;     //34pi/128
   sin[35]  =  14'b11001111100010;     //35pi/128
   cos[35]  =  14'b00101001110011;     //35pi/128
   sin[36]  =  14'b11001110100010;     //36pi/128
   cos[36]  =  14'b00101000100110;     //36pi/128
   sin[37]  =  14'b11001101100011;     //37pi/128
   cos[37]  =  14'b00100111010111;     //37pi/128
   sin[38]  =  14'b11001100100110;     //38pi/128
   cos[38]  =  14'b00100110000111;     //38pi/128
   sin[39]  =  14'b11001011101011;     //39pi/128
   cos[39]  =  14'b00100100110110;     //39pi/128
   sin[40]  =  14'b11001010110010;     //40pi/128
   cos[40]  =  14'b00100011100011;     //40pi/128
   sin[41]  =  14'b11001001111011;     //41pi/128
   cos[41]  =  14'b00100010001111;     //41pi/128
   sin[42]  =  14'b11001001000111;     //42pi/128
   cos[42]  =  14'b00100000111001;     //42pi/128
   sin[43]  =  14'b11001000010100;     //43pi/128
   cos[43]  =  14'b00011111100010;     //43pi/128
   sin[44]  =  14'b11000111100100;     //44pi/128
   cos[44]  =  14'b00011110001010;     //44pi/128
   sin[45]  =  14'b11000110110101;     //45pi/128
   cos[45]  =  14'b00011100110001;     //45pi/128
   sin[46]  =  14'b11000110001001;     //46pi/128
   cos[46]  =  14'b00011011010111;     //46pi/128
   sin[47]  =  14'b11000101011111;     //47pi/128
   cos[47]  =  14'b00011001111011;     //47pi/128
   sin[48]  =  14'b11000100111000;     //48pi/128
   cos[48]  =  14'b00011000011111;     //48pi/128
   sin[49]  =  14'b11000100010010;     //49pi/128
   cos[49]  =  14'b00010111000010;     //49pi/128
   sin[50]  =  14'b11000011101111;     //50pi/128
   cos[50]  =  14'b00010101100011;     //50pi/128
   sin[51]  =  14'b11000011001111;     //51pi/128
   cos[51]  =  14'b00010100000100;     //51pi/128
   sin[52]  =  14'b11000010110000;     //52pi/128
   cos[52]  =  14'b00010010100101;     //52pi/128
   sin[53]  =  14'b11000010010100;     //53pi/128
   cos[53]  =  14'b00010001000100;     //53pi/128
   sin[54]  =  14'b11000001111011;     //54pi/128
   cos[54]  =  14'b00001111100011;     //54pi/128
   sin[55]  =  14'b11000001100100;     //55pi/128
   cos[55]  =  14'b00001110000001;     //55pi/128
   sin[56]  =  14'b11000001001111;     //56pi/128
   cos[56]  =  14'b00001100011111;     //56pi/128
   sin[57]  =  14'b11000000111100;     //57pi/128
   cos[57]  =  14'b00001010111100;     //57pi/128
   sin[58]  =  14'b11000000101100;     //58pi/128
   cos[58]  =  14'b00001001011001;     //58pi/128
   sin[59]  =  14'b11000000011111;     //59pi/128
   cos[59]  =  14'b00000111110101;     //59pi/128
   sin[60]  =  14'b11000000010100;     //60pi/128
   cos[60]  =  14'b00000110010001;     //60pi/128
   sin[61]  =  14'b11000000001011;     //61pi/128
   cos[61]  =  14'b00000100101101;     //61pi/128
   sin[62]  =  14'b11000000000101;     //62pi/128
   cos[62]  =  14'b00000011001000;     //62pi/128
   sin[63]  =  14'b11000000000001;     //63pi/128
   cos[63]  =  14'b00000001100100;     //63pi/128
   sin[64]  =  14'b11000000000000;     //64pi/128
   cos[64]  =  14'b00000000000000;     //64pi/128
   sin[65]  =  14'b11000000000001;     //65pi/128
   cos[65]  =  14'b11111110011011;     //65pi/128
   sin[66]  =  14'b11000000000101;     //66pi/128
   cos[66]  =  14'b11111100110111;     //66pi/128
   sin[67]  =  14'b11000000001011;     //67pi/128
   cos[67]  =  14'b11111011010011;     //67pi/128
   sin[68]  =  14'b11000000010100;     //68pi/128
   cos[68]  =  14'b11111001101111;     //68pi/128
   sin[69]  =  14'b11000000011111;     //69pi/128
   cos[69]  =  14'b11111000001011;     //69pi/128
   sin[70]  =  14'b11000000101100;     //70pi/128
   cos[70]  =  14'b11110110100111;     //70pi/128
   sin[71]  =  14'b11000000111100;     //71pi/128
   cos[71]  =  14'b11110101000100;     //71pi/128
   sin[72]  =  14'b11000001001111;     //72pi/128
   cos[72]  =  14'b11110011100001;     //72pi/128
   sin[73]  =  14'b11000001100100;     //73pi/128
   cos[73]  =  14'b11110001111111;     //73pi/128
   sin[74]  =  14'b11000001111011;     //74pi/128
   cos[74]  =  14'b11110000011101;     //74pi/128
   sin[75]  =  14'b11000010010100;     //75pi/128
   cos[75]  =  14'b11101110111100;     //75pi/128
   sin[76]  =  14'b11000010110000;     //76pi/128
   cos[76]  =  14'b11101101011011;     //76pi/128
   sin[77]  =  14'b11000011001111;     //77pi/128
   cos[77]  =  14'b11101011111011;     //77pi/128
   sin[78]  =  14'b11000011101111;     //78pi/128
   cos[78]  =  14'b11101010011100;     //78pi/128
   sin[79]  =  14'b11000100010010;     //79pi/128
   cos[79]  =  14'b11101000111110;     //79pi/128
   sin[80]  =  14'b11000100111000;     //80pi/128
   cos[80]  =  14'b11100111100001;     //80pi/128
   sin[81]  =  14'b11000101011111;     //81pi/128
   cos[81]  =  14'b11100110000100;     //81pi/128
   sin[82]  =  14'b11000110001001;     //82pi/128
   cos[82]  =  14'b11100100101001;     //82pi/128
   sin[83]  =  14'b11000110110101;     //83pi/128
   cos[83]  =  14'b11100011001110;     //83pi/128
   sin[84]  =  14'b11000111100100;     //84pi/128
   cos[84]  =  14'b11100001110101;     //84pi/128
   sin[85]  =  14'b11001000010100;     //85pi/128
   cos[85]  =  14'b11100000011101;     //85pi/128
   sin[86]  =  14'b11001001000111;     //86pi/128
   cos[86]  =  14'b11011111000110;     //86pi/128
   sin[87]  =  14'b11001001111011;     //87pi/128
   cos[87]  =  14'b11011101110001;     //87pi/128
   sin[88]  =  14'b11001010110010;     //88pi/128
   cos[88]  =  14'b11011100011100;     //88pi/128
   sin[89]  =  14'b11001011101011;     //89pi/128
   cos[89]  =  14'b11011011001001;     //89pi/128
   sin[90]  =  14'b11001100100110;     //90pi/128
   cos[90]  =  14'b11011001111000;     //90pi/128
   sin[91]  =  14'b11001101100011;     //91pi/128
   cos[91]  =  14'b11011000101000;     //91pi/128
   sin[92]  =  14'b11001110100010;     //92pi/128
   cos[92]  =  14'b11010111011010;     //92pi/128
   sin[93]  =  14'b11001111100010;     //93pi/128
   cos[93]  =  14'b11010110001101;     //93pi/128
   sin[94]  =  14'b11010000100101;     //94pi/128
   cos[94]  =  14'b11010101000001;     //94pi/128
   sin[95]  =  14'b11010001101001;     //95pi/128
   cos[95]  =  14'b11010011111000;     //95pi/128
   sin[96]  =  14'b11010010110000;     //96pi/128
   cos[96]  =  14'b11010010110000;     //96pi/128
   sin[97]  =  14'b11010011111000;     //97pi/128
   cos[97]  =  14'b11010001101001;     //97pi/128
   sin[98]  =  14'b11010101000001;     //98pi/128
   cos[98]  =  14'b11010000100101;     //98pi/128
   sin[99]  =  14'b11010110001101;     //99pi/128
   cos[99]  =  14'b11001111100010;     //99pi/128
   sin[100]  =  14'b11010111011010;     //100pi/128
   cos[100]  =  14'b11001110100010;     //100pi/128
   sin[101]  =  14'b11011000101000;     //101pi/128
   cos[101]  =  14'b11001101100011;     //101pi/128
   sin[102]  =  14'b11011001111000;     //102pi/128
   cos[102]  =  14'b11001100100110;     //102pi/128
   sin[103]  =  14'b11011011001001;     //103pi/128
   cos[103]  =  14'b11001011101011;     //103pi/128
   sin[104]  =  14'b11011100011100;     //104pi/128
   cos[104]  =  14'b11001010110010;     //104pi/128
   sin[105]  =  14'b11011101110001;     //105pi/128
   cos[105]  =  14'b11001001111011;     //105pi/128
   sin[106]  =  14'b11011111000110;     //106pi/128
   cos[106]  =  14'b11001001000111;     //106pi/128
   sin[107]  =  14'b11100000011101;     //107pi/128
   cos[107]  =  14'b11001000010100;     //107pi/128
   sin[108]  =  14'b11100001110101;     //108pi/128
   cos[108]  =  14'b11000111100100;     //108pi/128
   sin[109]  =  14'b11100011001110;     //109pi/128
   cos[109]  =  14'b11000110110101;     //109pi/128
   sin[110]  =  14'b11100100101001;     //110pi/128
   cos[110]  =  14'b11000110001001;     //110pi/128
   sin[111]  =  14'b11100110000100;     //111pi/128
   cos[111]  =  14'b11000101011111;     //111pi/128
   sin[112]  =  14'b11100111100001;     //112pi/128
   cos[112]  =  14'b11000100111000;     //112pi/128
   sin[113]  =  14'b11101000111110;     //113pi/128
   cos[113]  =  14'b11000100010010;     //113pi/128
   sin[114]  =  14'b11101010011100;     //114pi/128
   cos[114]  =  14'b11000011101111;     //114pi/128
   sin[115]  =  14'b11101011111011;     //115pi/128
   cos[115]  =  14'b11000011001111;     //115pi/128
   sin[116]  =  14'b11101101011011;     //116pi/128
   cos[116]  =  14'b11000010110000;     //116pi/128
   sin[117]  =  14'b11101110111100;     //117pi/128
   cos[117]  =  14'b11000010010100;     //117pi/128
   sin[118]  =  14'b11110000011101;     //118pi/128
   cos[118]  =  14'b11000001111011;     //118pi/128
   sin[119]  =  14'b11110001111111;     //119pi/128
   cos[119]  =  14'b11000001100100;     //119pi/128
   sin[120]  =  14'b11110011100001;     //120pi/128
   cos[120]  =  14'b11000001001111;     //120pi/128
   sin[121]  =  14'b11110101000100;     //121pi/128
   cos[121]  =  14'b11000000111100;     //121pi/128
   sin[122]  =  14'b11110110100111;     //122pi/128
   cos[122]  =  14'b11000000101100;     //122pi/128
   sin[123]  =  14'b11111000001011;     //123pi/128
   cos[123]  =  14'b11000000011111;     //123pi/128
   sin[124]  =  14'b11111001101111;     //124pi/128
   cos[124]  =  14'b11000000010100;     //124pi/128
   sin[125]  =  14'b11111011010011;     //125pi/128
   cos[125]  =  14'b11000000001011;     //125pi/128
   sin[126]  =  14'b11111100110111;     //126pi/128
   cos[126]  =  14'b11000000000101;     //126pi/128
   sin[127]  =  14'b11111110011011;     //127pi/128
   cos[127]  =  14'b11000000000001;     //127pi/128

   sin[128]  =  14'b00000000000000;     //0pi/128
   cos[128]  =  14'b01000000000000;     //0pi/128
   sin[129]  =  14'b11111110110000;     //1pi/128
   cos[129]  =  14'b00111111111111;     //1pi/128
   sin[130]  =  14'b11111101011111;     //2pi/128
   cos[130]  =  14'b00111111111100;     //2pi/128
   sin[131]  =  14'b11111100001111;     //3pi/128
   cos[131]  =  14'b00111111111000;     //3pi/128
   sin[132]  =  14'b11111010111111;     //4pi/128
   cos[132]  =  14'b00111111110011;     //4pi/128
   sin[133]  =  14'b11111001101111;     //5pi/128
   cos[133]  =  14'b00111111101100;     //5pi/128
   sin[134]  =  14'b11111000011111;     //6pi/128
   cos[134]  =  14'b00111111100011;     //6pi/128
   sin[135]  =  14'b11110111001111;     //7pi/128
   cos[135]  =  14'b00111111011001;     //7pi/128
   sin[136]  =  14'b11110101111111;     //8pi/128
   cos[136]  =  14'b00111111001101;     //8pi/128
   sin[137]  =  14'b11110100110000;     //9pi/128
   cos[137]  =  14'b00111111000000;     //9pi/128
   sin[138]  =  14'b11110011100001;     //10pi/128
   cos[138]  =  14'b00111110110001;     //10pi/128
   sin[139]  =  14'b11110010010010;     //11pi/128
   cos[139]  =  14'b00111110100000;     //11pi/128
   sin[140]  =  14'b11110001000100;     //12pi/128
   cos[140]  =  14'b00111110001110;     //12pi/128
   sin[141]  =  14'b11101111110110;     //13pi/128
   cos[141]  =  14'b00111101111011;     //13pi/128
   sin[142]  =  14'b11101110101000;     //14pi/128
   cos[142]  =  14'b00111101100110;     //14pi/128
   sin[143]  =  14'b11101101011011;     //15pi/128
   cos[143]  =  14'b00111101001111;     //15pi/128
   sin[144]  =  14'b11101100001110;     //16pi/128
   cos[144]  =  14'b00111100110111;     //16pi/128
   sin[145]  =  14'b11101011000010;     //17pi/128
   cos[145]  =  14'b00111100011101;     //17pi/128
   sin[146]  =  14'b11101001110110;     //18pi/128
   cos[146]  =  14'b00111100000010;     //18pi/128
   sin[147]  =  14'b11101000101011;     //19pi/128
   cos[147]  =  14'b00111011100110;     //19pi/128
   sin[148]  =  14'b11100111100001;     //20pi/128
   cos[148]  =  14'b00111011001000;     //20pi/128
   sin[149]  =  14'b11100110010111;     //21pi/128
   cos[149]  =  14'b00111010101000;     //21pi/128
   sin[150]  =  14'b11100101001101;     //22pi/128
   cos[150]  =  14'b00111010000111;     //22pi/128
   sin[151]  =  14'b11100100000100;     //23pi/128
   cos[151]  =  14'b00111001100101;     //23pi/128
   sin[152]  =  14'b11100010111100;     //24pi/128
   cos[152]  =  14'b00111001000001;     //24pi/128
   sin[153]  =  14'b11100001110101;     //25pi/128
   cos[153]  =  14'b00111000011100;     //25pi/128
   sin[154]  =  14'b11100000101111;     //26pi/128
   cos[154]  =  14'b00110111110101;     //26pi/128
   sin[155]  =  14'b11011111101001;     //27pi/128
   cos[155]  =  14'b00110111001101;     //27pi/128
   sin[156]  =  14'b11011110100100;     //28pi/128
   cos[156]  =  14'b00110110100100;     //28pi/128
   sin[157]  =  14'b11011101100000;     //29pi/128
   cos[157]  =  14'b00110101111001;     //29pi/128
   sin[158]  =  14'b11011100011100;     //30pi/128
   cos[158]  =  14'b00110101001101;     //30pi/128
   sin[159]  =  14'b11011011011010;     //31pi/128
   cos[159]  =  14'b00110100100000;     //31pi/128
   sin[160]  =  14'b11011010011000;     //32pi/128
   cos[160]  =  14'b00110011110001;     //32pi/128
   sin[161]  =  14'b11011001011000;     //33pi/128
   cos[161]  =  14'b00110011000001;     //33pi/128
   sin[162]  =  14'b11011000011000;     //34pi/128
   cos[162]  =  14'b00110010010000;     //34pi/128
   sin[163]  =  14'b11010111011010;     //35pi/128
   cos[163]  =  14'b00110001011110;     //35pi/128
   sin[164]  =  14'b11010110011100;     //36pi/128
   cos[164]  =  14'b00110000101010;     //36pi/128
   sin[165]  =  14'b11010101011111;     //37pi/128
   cos[165]  =  14'b00101111110101;     //37pi/128
   sin[166]  =  14'b11010100100100;     //38pi/128
   cos[166]  =  14'b00101110111111;     //38pi/128
   sin[167]  =  14'b11010011101001;     //39pi/128
   cos[167]  =  14'b00101110001000;     //39pi/128
   sin[168]  =  14'b11010010110000;     //40pi/128
   cos[168]  =  14'b00101101010000;     //40pi/128
   sin[169]  =  14'b11010001110111;     //41pi/128
   cos[169]  =  14'b00101100010110;     //41pi/128
   sin[170]  =  14'b11010001000000;     //42pi/128
   cos[170]  =  14'b00101011011100;     //42pi/128
   sin[171]  =  14'b11010000001010;     //43pi/128
   cos[171]  =  14'b00101010100000;     //43pi/128
   sin[172]  =  14'b11001111010101;     //44pi/128
   cos[172]  =  14'b00101001100100;     //44pi/128
   sin[173]  =  14'b11001110100010;     //45pi/128
   cos[173]  =  14'b00101000100110;     //45pi/128
   sin[174]  =  14'b11001101101111;     //46pi/128
   cos[174]  =  14'b00100111100111;     //46pi/128
   sin[175]  =  14'b11001100111110;     //47pi/128
   cos[175]  =  14'b00100110101000;     //47pi/128
   sin[176]  =  14'b11001100001110;     //48pi/128
   cos[176]  =  14'b00100101100111;     //48pi/128
   sin[177]  =  14'b11001011100000;     //49pi/128
   cos[177]  =  14'b00100100100110;     //49pi/128
   sin[178]  =  14'b11001010110010;     //50pi/128
   cos[178]  =  14'b00100011100011;     //50pi/128
   sin[179]  =  14'b11001010000110;     //51pi/128
   cos[179]  =  14'b00100010100000;     //51pi/128
   sin[180]  =  14'b11001001011100;     //52pi/128
   cos[180]  =  14'b00100001011100;     //52pi/128
   sin[181]  =  14'b11001000110010;     //53pi/128
   cos[181]  =  14'b00100000010111;     //53pi/128
   sin[182]  =  14'b11001000001010;     //54pi/128
   cos[182]  =  14'b00011111010001;     //54pi/128
   sin[183]  =  14'b11000111100100;     //55pi/128
   cos[183]  =  14'b00011110001010;     //55pi/128
   sin[184]  =  14'b11000110111110;     //56pi/128
   cos[184]  =  14'b00011101000011;     //56pi/128
   sin[185]  =  14'b11000110011011;     //57pi/128
   cos[185]  =  14'b00011011111011;     //57pi/128
   sin[186]  =  14'b11000101111000;     //58pi/128
   cos[186]  =  14'b00011010110010;     //58pi/128
   sin[187]  =  14'b11000101010111;     //59pi/128
   cos[187]  =  14'b00011001101001;     //59pi/128
   sin[188]  =  14'b11000100111000;     //60pi/128
   cos[188]  =  14'b00011000011111;     //60pi/128
   sin[189]  =  14'b11000100011010;     //61pi/128
   cos[189]  =  14'b00010111010100;     //61pi/128
   sin[190]  =  14'b11000011111101;     //62pi/128
   cos[190]  =  14'b00010110001001;     //62pi/128
   sin[191]  =  14'b11000011100010;     //63pi/128
   cos[191]  =  14'b00010100111101;     //63pi/128
   sin[192]  =  14'b11000011001000;     //64pi/128
   cos[192]  =  14'b00010011110001;     //64pi/128
   sin[193]  =  14'b11000010110000;     //65pi/128
   cos[193]  =  14'b00010010100101;     //65pi/128
   sin[194]  =  14'b11000010011010;     //66pi/128
   cos[194]  =  14'b00010001010111;     //66pi/128
   sin[195]  =  14'b11000010000101;     //67pi/128
   cos[195]  =  14'b00010000001010;     //67pi/128
   sin[196]  =  14'b11000001110001;     //68pi/128
   cos[196]  =  14'b00001110111100;     //68pi/128
   sin[197]  =  14'b11000001011111;     //69pi/128
   cos[197]  =  14'b00001101101101;     //69pi/128
   sin[198]  =  14'b11000001001111;     //70pi/128
   cos[198]  =  14'b00001100011111;     //70pi/128
   sin[199]  =  14'b11000001000000;     //71pi/128
   cos[199]  =  14'b00001011010000;     //71pi/128
   sin[200]  =  14'b11000000110010;     //72pi/128
   cos[200]  =  14'b00001010000000;     //72pi/128
   sin[201]  =  14'b11000000100111;     //73pi/128
   cos[201]  =  14'b00001000110001;     //73pi/128
   sin[202]  =  14'b11000000011100;     //74pi/128
   cos[202]  =  14'b00000111100001;     //74pi/128
   sin[203]  =  14'b11000000010100;     //75pi/128
   cos[203]  =  14'b00000110010001;     //75pi/128
   sin[204]  =  14'b11000000001101;     //76pi/128
   cos[204]  =  14'b00000101000001;     //76pi/128
   sin[205]  =  14'b11000000000111;     //77pi/128
   cos[205]  =  14'b00000011110001;     //77pi/128
   sin[206]  =  14'b11000000000011;     //78pi/128
   cos[206]  =  14'b00000010100000;     //78pi/128
   sin[207]  =  14'b11000000000001;     //79pi/128
   cos[207]  =  14'b00000001010000;     //79pi/128
   sin[208]  =  14'b11000000000000;     //80pi/128
   cos[208]  =  14'b00000000000000;     //80pi/128
   sin[209]  =  14'b11000000000001;     //81pi/128
   cos[209]  =  14'b11111110110000;     //81pi/128
   sin[210]  =  14'b11000000000011;     //82pi/128
   cos[210]  =  14'b11111101011111;     //82pi/128
   sin[211]  =  14'b11000000000111;     //83pi/128
   cos[211]  =  14'b11111100001111;     //83pi/128
   sin[212]  =  14'b11000000001101;     //84pi/128
   cos[212]  =  14'b11111010111111;     //84pi/128
   sin[213]  =  14'b11000000010100;     //85pi/128
   cos[213]  =  14'b11111001101111;     //85pi/128
   sin[214]  =  14'b11000000011100;     //86pi/128
   cos[214]  =  14'b11111000011111;     //86pi/128
   sin[215]  =  14'b11000000100111;     //87pi/128
   cos[215]  =  14'b11110111001111;     //87pi/128
   sin[216]  =  14'b11000000110010;     //88pi/128
   cos[216]  =  14'b11110101111111;     //88pi/128
   sin[217]  =  14'b11000001000000;     //89pi/128
   cos[217]  =  14'b11110100110000;     //89pi/128
   sin[218]  =  14'b11000001001111;     //90pi/128
   cos[218]  =  14'b11110011100001;     //90pi/128
   sin[219]  =  14'b11000001011111;     //91pi/128
   cos[219]  =  14'b11110010010010;     //91pi/128
   sin[220]  =  14'b11000001110001;     //92pi/128
   cos[220]  =  14'b11110001000100;     //92pi/128
   sin[221]  =  14'b11000010000101;     //93pi/128
   cos[221]  =  14'b11101111110110;     //93pi/128
   sin[222]  =  14'b11000010011010;     //94pi/128
   cos[222]  =  14'b11101110101000;     //94pi/128
   sin[223]  =  14'b11000010110000;     //95pi/128
   cos[223]  =  14'b11101101011011;     //95pi/128
   sin[224]  =  14'b11000011001000;     //96pi/128
   cos[224]  =  14'b11101100001110;     //96pi/128
   sin[225]  =  14'b11000011100010;     //97pi/128
   cos[225]  =  14'b11101011000010;     //97pi/128
   sin[226]  =  14'b11000011111101;     //98pi/128
   cos[226]  =  14'b11101001110110;     //98pi/128
   sin[227]  =  14'b11000100011010;     //99pi/128
   cos[227]  =  14'b11101000101011;     //99pi/128
   sin[228]  =  14'b11000100111000;     //100pi/128
   cos[228]  =  14'b11100111100001;     //100pi/128
   sin[229]  =  14'b11000101010111;     //101pi/128
   cos[229]  =  14'b11100110010111;     //101pi/128
   sin[230]  =  14'b11000101111000;     //102pi/128
   cos[230]  =  14'b11100101001101;     //102pi/128
   sin[231]  =  14'b11000110011011;     //103pi/128
   cos[231]  =  14'b11100100000100;     //103pi/128
   sin[232]  =  14'b11000110111110;     //104pi/128
   cos[232]  =  14'b11100010111100;     //104pi/128
   sin[233]  =  14'b11000111100100;     //105pi/128
   cos[233]  =  14'b11100001110101;     //105pi/128
   sin[234]  =  14'b11001000001010;     //106pi/128
   cos[234]  =  14'b11100000101111;     //106pi/128
   sin[235]  =  14'b11001000110010;     //107pi/128
   cos[235]  =  14'b11011111101001;     //107pi/128
   sin[236]  =  14'b11001001011100;     //108pi/128
   cos[236]  =  14'b11011110100100;     //108pi/128
   sin[237]  =  14'b11001010000110;     //109pi/128
   cos[237]  =  14'b11011101100000;     //109pi/128
   sin[238]  =  14'b11001010110010;     //110pi/128
   cos[238]  =  14'b11011100011100;     //110pi/128
   sin[239]  =  14'b11001011100000;     //111pi/128
   cos[239]  =  14'b11011011011010;     //111pi/128
   sin[240]  =  14'b11001100001110;     //112pi/128
   cos[240]  =  14'b11011010011000;     //112pi/128
   sin[241]  =  14'b11001100111110;     //113pi/128
   cos[241]  =  14'b11011001011000;     //113pi/128
   sin[242]  =  14'b11001101101111;     //114pi/128
   cos[242]  =  14'b11011000011000;     //114pi/128
   sin[243]  =  14'b11001110100010;     //115pi/128
   cos[243]  =  14'b11010111011010;     //115pi/128
   sin[244]  =  14'b11001111010101;     //116pi/128
   cos[244]  =  14'b11010110011100;     //116pi/128
   sin[245]  =  14'b11010000001010;     //117pi/128
   cos[245]  =  14'b11010101011111;     //117pi/128
   sin[246]  =  14'b11010001000000;     //118pi/128
   cos[246]  =  14'b11010100100100;     //118pi/128
   sin[247]  =  14'b11010001110111;     //119pi/128
   cos[247]  =  14'b11010011101001;     //119pi/128
   sin[248]  =  14'b11010010110000;     //120pi/128
   cos[248]  =  14'b11010010110000;     //120pi/128
   sin[249]  =  14'b11010011101001;     //121pi/128
   cos[249]  =  14'b11010001110111;     //121pi/128
   sin[250]  =  14'b11010100100100;     //122pi/128
   cos[250]  =  14'b11010001000000;     //122pi/128
   sin[251]  =  14'b11010101011111;     //123pi/128
   cos[251]  =  14'b11010000001010;     //123pi/128
   sin[252]  =  14'b11010110011100;     //124pi/128
   cos[252]  =  14'b11001111010101;     //124pi/128
   sin[253]  =  14'b11010111011010;     //125pi/128
   cos[253]  =  14'b11001110100010;     //125pi/128
   sin[254]  =  14'b11011000011000;     //126pi/128
   cos[254]  =  14'b11001101101111;     //126pi/128
   sin[255]  =  14'b11011001011000;     //127pi/128
   cos[255]  =  14'b11001100111110;     //127pi/128
end
endmodule