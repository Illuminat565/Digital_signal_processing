module  M_TWIDLE_6_bit #(parameter SIZE =10, word_length_tw = 6) (
    input            clk,
    input            en_rd, 
    input   [10:0]   rd_ptr_angle,
    input            en_modf, 

    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );


reg signed [word_length_tw-1:0]  cos  [511:0];
reg signed [word_length_tw-1:0]  sin  [511:0];

reg signed [word_length_tw-1:0]  m_cos  [511:0];
reg signed [word_length_tw-1:0]  m_sin  [511:0];

reg signed [word_length_tw-1:0]  cos_temp;
reg signed [word_length_tw-1:0]  sin_temp;

reg signed [word_length_tw-1:0]  m_cos_temp;
reg signed [word_length_tw-1:0]  m_sin_temp;


//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & ~ en_modf ) begin
                  cos_temp           <= cos   [rd_ptr_angle];
                  sin_temp           <= sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd & en_modf ) begin
                  m_cos_temp           <= m_cos   [rd_ptr_angle];
                  m_sin_temp           <= m_sin   [rd_ptr_angle];
             end 
        end
//--------------------------------handle read tw factor------------------------------
     always @(*) begin 
             if (en_modf ) begin
                  cos_data           <= m_cos_temp;
                  sin_data           <= m_sin_temp;
             end else begin
                  cos_data           <= cos_temp;
                  sin_data           <= sin_temp;
             end
        end
//----------------------------------------------------------------------------------------
initial begin

   sin[0]  =  6'b000000;     //0pi/512
   cos[0]  =  6'b010000;     //0pi/512
   sin[1]  =  6'b000000;     //1pi/512
   cos[1]  =  6'b001111;     //1pi/512
   sin[2]  =  6'b000000;     //2pi/512
   cos[2]  =  6'b001111;     //2pi/512
   sin[3]  =  6'b000000;     //3pi/512
   cos[3]  =  6'b001111;     //3pi/512
   sin[4]  =  6'b000000;     //4pi/512
   cos[4]  =  6'b001111;     //4pi/512
   sin[5]  =  6'b000000;     //5pi/512
   cos[5]  =  6'b001111;     //5pi/512
   sin[6]  =  6'b111111;     //6pi/512
   cos[6]  =  6'b001111;     //6pi/512
   sin[7]  =  6'b111111;     //7pi/512
   cos[7]  =  6'b001111;     //7pi/512
   sin[8]  =  6'b111111;     //8pi/512
   cos[8]  =  6'b001111;     //8pi/512
   sin[9]  =  6'b111111;     //9pi/512
   cos[9]  =  6'b001111;     //9pi/512
   sin[10]  =  6'b111111;     //10pi/512
   cos[10]  =  6'b001111;     //10pi/512
   sin[11]  =  6'b111111;     //11pi/512
   cos[11]  =  6'b001111;     //11pi/512
   sin[12]  =  6'b111111;     //12pi/512
   cos[12]  =  6'b001111;     //12pi/512
   sin[13]  =  6'b111111;     //13pi/512
   cos[13]  =  6'b001111;     //13pi/512
   sin[14]  =  6'b111111;     //14pi/512
   cos[14]  =  6'b001111;     //14pi/512
   sin[15]  =  6'b111111;     //15pi/512
   cos[15]  =  6'b001111;     //15pi/512
   sin[16]  =  6'b111110;     //16pi/512
   cos[16]  =  6'b001111;     //16pi/512
   sin[17]  =  6'b111110;     //17pi/512
   cos[17]  =  6'b001111;     //17pi/512
   sin[18]  =  6'b111110;     //18pi/512
   cos[18]  =  6'b001111;     //18pi/512
   sin[19]  =  6'b111110;     //19pi/512
   cos[19]  =  6'b001111;     //19pi/512
   sin[20]  =  6'b111110;     //20pi/512
   cos[20]  =  6'b001111;     //20pi/512
   sin[21]  =  6'b111110;     //21pi/512
   cos[21]  =  6'b001111;     //21pi/512
   sin[22]  =  6'b111110;     //22pi/512
   cos[22]  =  6'b001111;     //22pi/512
   sin[23]  =  6'b111110;     //23pi/512
   cos[23]  =  6'b001111;     //23pi/512
   sin[24]  =  6'b111110;     //24pi/512
   cos[24]  =  6'b001111;     //24pi/512
   sin[25]  =  6'b111110;     //25pi/512
   cos[25]  =  6'b001111;     //25pi/512
   sin[26]  =  6'b111101;     //26pi/512
   cos[26]  =  6'b001111;     //26pi/512
   sin[27]  =  6'b111101;     //27pi/512
   cos[27]  =  6'b001111;     //27pi/512
   sin[28]  =  6'b111101;     //28pi/512
   cos[28]  =  6'b001111;     //28pi/512
   sin[29]  =  6'b111101;     //29pi/512
   cos[29]  =  6'b001111;     //29pi/512
   sin[30]  =  6'b111101;     //30pi/512
   cos[30]  =  6'b001111;     //30pi/512
   sin[31]  =  6'b111101;     //31pi/512
   cos[31]  =  6'b001111;     //31pi/512
   sin[32]  =  6'b111101;     //32pi/512
   cos[32]  =  6'b001111;     //32pi/512
   sin[33]  =  6'b111101;     //33pi/512
   cos[33]  =  6'b001111;     //33pi/512
   sin[34]  =  6'b111101;     //34pi/512
   cos[34]  =  6'b001111;     //34pi/512
   sin[35]  =  6'b111101;     //35pi/512
   cos[35]  =  6'b001111;     //35pi/512
   sin[36]  =  6'b111100;     //36pi/512
   cos[36]  =  6'b001111;     //36pi/512
   sin[37]  =  6'b111100;     //37pi/512
   cos[37]  =  6'b001111;     //37pi/512
   sin[38]  =  6'b111100;     //38pi/512
   cos[38]  =  6'b001111;     //38pi/512
   sin[39]  =  6'b111100;     //39pi/512
   cos[39]  =  6'b001111;     //39pi/512
   sin[40]  =  6'b111100;     //40pi/512
   cos[40]  =  6'b001111;     //40pi/512
   sin[41]  =  6'b111100;     //41pi/512
   cos[41]  =  6'b001111;     //41pi/512
   sin[42]  =  6'b111100;     //42pi/512
   cos[42]  =  6'b001111;     //42pi/512
   sin[43]  =  6'b111100;     //43pi/512
   cos[43]  =  6'b001111;     //43pi/512
   sin[44]  =  6'b111100;     //44pi/512
   cos[44]  =  6'b001111;     //44pi/512
   sin[45]  =  6'b111100;     //45pi/512
   cos[45]  =  6'b001111;     //45pi/512
   sin[46]  =  6'b111100;     //46pi/512
   cos[46]  =  6'b001111;     //46pi/512
   sin[47]  =  6'b111011;     //47pi/512
   cos[47]  =  6'b001111;     //47pi/512
   sin[48]  =  6'b111011;     //48pi/512
   cos[48]  =  6'b001111;     //48pi/512
   sin[49]  =  6'b111011;     //49pi/512
   cos[49]  =  6'b001111;     //49pi/512
   sin[50]  =  6'b111011;     //50pi/512
   cos[50]  =  6'b001111;     //50pi/512
   sin[51]  =  6'b111011;     //51pi/512
   cos[51]  =  6'b001111;     //51pi/512
   sin[52]  =  6'b111011;     //52pi/512
   cos[52]  =  6'b001111;     //52pi/512
   sin[53]  =  6'b111011;     //53pi/512
   cos[53]  =  6'b001111;     //53pi/512
   sin[54]  =  6'b111011;     //54pi/512
   cos[54]  =  6'b001111;     //54pi/512
   sin[55]  =  6'b111011;     //55pi/512
   cos[55]  =  6'b001111;     //55pi/512
   sin[56]  =  6'b111011;     //56pi/512
   cos[56]  =  6'b001111;     //56pi/512
   sin[57]  =  6'b111011;     //57pi/512
   cos[57]  =  6'b001111;     //57pi/512
   sin[58]  =  6'b111010;     //58pi/512
   cos[58]  =  6'b001110;     //58pi/512
   sin[59]  =  6'b111010;     //59pi/512
   cos[59]  =  6'b001110;     //59pi/512
   sin[60]  =  6'b111010;     //60pi/512
   cos[60]  =  6'b001110;     //60pi/512
   sin[61]  =  6'b111010;     //61pi/512
   cos[61]  =  6'b001110;     //61pi/512
   sin[62]  =  6'b111010;     //62pi/512
   cos[62]  =  6'b001110;     //62pi/512
   sin[63]  =  6'b111010;     //63pi/512
   cos[63]  =  6'b001110;     //63pi/512
   sin[64]  =  6'b111010;     //64pi/512
   cos[64]  =  6'b001110;     //64pi/512
   sin[65]  =  6'b111010;     //65pi/512
   cos[65]  =  6'b001110;     //65pi/512
   sin[66]  =  6'b111010;     //66pi/512
   cos[66]  =  6'b001110;     //66pi/512
   sin[67]  =  6'b111010;     //67pi/512
   cos[67]  =  6'b001110;     //67pi/512
   sin[68]  =  6'b111010;     //68pi/512
   cos[68]  =  6'b001110;     //68pi/512
   sin[69]  =  6'b111001;     //69pi/512
   cos[69]  =  6'b001110;     //69pi/512
   sin[70]  =  6'b111001;     //70pi/512
   cos[70]  =  6'b001110;     //70pi/512
   sin[71]  =  6'b111001;     //71pi/512
   cos[71]  =  6'b001110;     //71pi/512
   sin[72]  =  6'b111001;     //72pi/512
   cos[72]  =  6'b001110;     //72pi/512
   sin[73]  =  6'b111001;     //73pi/512
   cos[73]  =  6'b001110;     //73pi/512
   sin[74]  =  6'b111001;     //74pi/512
   cos[74]  =  6'b001110;     //74pi/512
   sin[75]  =  6'b111001;     //75pi/512
   cos[75]  =  6'b001110;     //75pi/512
   sin[76]  =  6'b111001;     //76pi/512
   cos[76]  =  6'b001110;     //76pi/512
   sin[77]  =  6'b111001;     //77pi/512
   cos[77]  =  6'b001110;     //77pi/512
   sin[78]  =  6'b111001;     //78pi/512
   cos[78]  =  6'b001110;     //78pi/512
   sin[79]  =  6'b111001;     //79pi/512
   cos[79]  =  6'b001110;     //79pi/512
   sin[80]  =  6'b111000;     //80pi/512
   cos[80]  =  6'b001110;     //80pi/512
   sin[81]  =  6'b111000;     //81pi/512
   cos[81]  =  6'b001110;     //81pi/512
   sin[82]  =  6'b111000;     //82pi/512
   cos[82]  =  6'b001110;     //82pi/512
   sin[83]  =  6'b111000;     //83pi/512
   cos[83]  =  6'b001101;     //83pi/512
   sin[84]  =  6'b111000;     //84pi/512
   cos[84]  =  6'b001101;     //84pi/512
   sin[85]  =  6'b111000;     //85pi/512
   cos[85]  =  6'b001101;     //85pi/512
   sin[86]  =  6'b111000;     //86pi/512
   cos[86]  =  6'b001101;     //86pi/512
   sin[87]  =  6'b111000;     //87pi/512
   cos[87]  =  6'b001101;     //87pi/512
   sin[88]  =  6'b111000;     //88pi/512
   cos[88]  =  6'b001101;     //88pi/512
   sin[89]  =  6'b111000;     //89pi/512
   cos[89]  =  6'b001101;     //89pi/512
   sin[90]  =  6'b111000;     //90pi/512
   cos[90]  =  6'b001101;     //90pi/512
   sin[91]  =  6'b111000;     //91pi/512
   cos[91]  =  6'b001101;     //91pi/512
   sin[92]  =  6'b110111;     //92pi/512
   cos[92]  =  6'b001101;     //92pi/512
   sin[93]  =  6'b110111;     //93pi/512
   cos[93]  =  6'b001101;     //93pi/512
   sin[94]  =  6'b110111;     //94pi/512
   cos[94]  =  6'b001101;     //94pi/512
   sin[95]  =  6'b110111;     //95pi/512
   cos[95]  =  6'b001101;     //95pi/512
   sin[96]  =  6'b110111;     //96pi/512
   cos[96]  =  6'b001101;     //96pi/512
   sin[97]  =  6'b110111;     //97pi/512
   cos[97]  =  6'b001101;     //97pi/512
   sin[98]  =  6'b110111;     //98pi/512
   cos[98]  =  6'b001101;     //98pi/512
   sin[99]  =  6'b110111;     //99pi/512
   cos[99]  =  6'b001101;     //99pi/512
   sin[100]  =  6'b110111;     //100pi/512
   cos[100]  =  6'b001101;     //100pi/512
   sin[101]  =  6'b110111;     //101pi/512
   cos[101]  =  6'b001101;     //101pi/512
   sin[102]  =  6'b110111;     //102pi/512
   cos[102]  =  6'b001100;     //102pi/512
   sin[103]  =  6'b110111;     //103pi/512
   cos[103]  =  6'b001100;     //103pi/512
   sin[104]  =  6'b110110;     //104pi/512
   cos[104]  =  6'b001100;     //104pi/512
   sin[105]  =  6'b110110;     //105pi/512
   cos[105]  =  6'b001100;     //105pi/512
   sin[106]  =  6'b110110;     //106pi/512
   cos[106]  =  6'b001100;     //106pi/512
   sin[107]  =  6'b110110;     //107pi/512
   cos[107]  =  6'b001100;     //107pi/512
   sin[108]  =  6'b110110;     //108pi/512
   cos[108]  =  6'b001100;     //108pi/512
   sin[109]  =  6'b110110;     //109pi/512
   cos[109]  =  6'b001100;     //109pi/512
   sin[110]  =  6'b110110;     //110pi/512
   cos[110]  =  6'b001100;     //110pi/512
   sin[111]  =  6'b110110;     //111pi/512
   cos[111]  =  6'b001100;     //111pi/512
   sin[112]  =  6'b110110;     //112pi/512
   cos[112]  =  6'b001100;     //112pi/512
   sin[113]  =  6'b110110;     //113pi/512
   cos[113]  =  6'b001100;     //113pi/512
   sin[114]  =  6'b110110;     //114pi/512
   cos[114]  =  6'b001100;     //114pi/512
   sin[115]  =  6'b110110;     //115pi/512
   cos[115]  =  6'b001100;     //115pi/512
   sin[116]  =  6'b110110;     //116pi/512
   cos[116]  =  6'b001100;     //116pi/512
   sin[117]  =  6'b110101;     //117pi/512
   cos[117]  =  6'b001100;     //117pi/512
   sin[118]  =  6'b110101;     //118pi/512
   cos[118]  =  6'b001011;     //118pi/512
   sin[119]  =  6'b110101;     //119pi/512
   cos[119]  =  6'b001011;     //119pi/512
   sin[120]  =  6'b110101;     //120pi/512
   cos[120]  =  6'b001011;     //120pi/512
   sin[121]  =  6'b110101;     //121pi/512
   cos[121]  =  6'b001011;     //121pi/512
   sin[122]  =  6'b110101;     //122pi/512
   cos[122]  =  6'b001011;     //122pi/512
   sin[123]  =  6'b110101;     //123pi/512
   cos[123]  =  6'b001011;     //123pi/512
   sin[124]  =  6'b110101;     //124pi/512
   cos[124]  =  6'b001011;     //124pi/512
   sin[125]  =  6'b110101;     //125pi/512
   cos[125]  =  6'b001011;     //125pi/512
   sin[126]  =  6'b110101;     //126pi/512
   cos[126]  =  6'b001011;     //126pi/512
   sin[127]  =  6'b110101;     //127pi/512
   cos[127]  =  6'b001011;     //127pi/512
   sin[128]  =  6'b110101;     //128pi/512
   cos[128]  =  6'b001011;     //128pi/512
   sin[129]  =  6'b110101;     //129pi/512
   cos[129]  =  6'b001011;     //129pi/512
   sin[130]  =  6'b110101;     //130pi/512
   cos[130]  =  6'b001011;     //130pi/512
   sin[131]  =  6'b110100;     //131pi/512
   cos[131]  =  6'b001011;     //131pi/512
   sin[132]  =  6'b110100;     //132pi/512
   cos[132]  =  6'b001011;     //132pi/512
   sin[133]  =  6'b110100;     //133pi/512
   cos[133]  =  6'b001010;     //133pi/512
   sin[134]  =  6'b110100;     //134pi/512
   cos[134]  =  6'b001010;     //134pi/512
   sin[135]  =  6'b110100;     //135pi/512
   cos[135]  =  6'b001010;     //135pi/512
   sin[136]  =  6'b110100;     //136pi/512
   cos[136]  =  6'b001010;     //136pi/512
   sin[137]  =  6'b110100;     //137pi/512
   cos[137]  =  6'b001010;     //137pi/512
   sin[138]  =  6'b110100;     //138pi/512
   cos[138]  =  6'b001010;     //138pi/512
   sin[139]  =  6'b110100;     //139pi/512
   cos[139]  =  6'b001010;     //139pi/512
   sin[140]  =  6'b110100;     //140pi/512
   cos[140]  =  6'b001010;     //140pi/512
   sin[141]  =  6'b110100;     //141pi/512
   cos[141]  =  6'b001010;     //141pi/512
   sin[142]  =  6'b110100;     //142pi/512
   cos[142]  =  6'b001010;     //142pi/512
   sin[143]  =  6'b110100;     //143pi/512
   cos[143]  =  6'b001010;     //143pi/512
   sin[144]  =  6'b110100;     //144pi/512
   cos[144]  =  6'b001010;     //144pi/512
   sin[145]  =  6'b110100;     //145pi/512
   cos[145]  =  6'b001010;     //145pi/512
   sin[146]  =  6'b110100;     //146pi/512
   cos[146]  =  6'b001001;     //146pi/512
   sin[147]  =  6'b110011;     //147pi/512
   cos[147]  =  6'b001001;     //147pi/512
   sin[148]  =  6'b110011;     //148pi/512
   cos[148]  =  6'b001001;     //148pi/512
   sin[149]  =  6'b110011;     //149pi/512
   cos[149]  =  6'b001001;     //149pi/512
   sin[150]  =  6'b110011;     //150pi/512
   cos[150]  =  6'b001001;     //150pi/512
   sin[151]  =  6'b110011;     //151pi/512
   cos[151]  =  6'b001001;     //151pi/512
   sin[152]  =  6'b110011;     //152pi/512
   cos[152]  =  6'b001001;     //152pi/512
   sin[153]  =  6'b110011;     //153pi/512
   cos[153]  =  6'b001001;     //153pi/512
   sin[154]  =  6'b110011;     //154pi/512
   cos[154]  =  6'b001001;     //154pi/512
   sin[155]  =  6'b110011;     //155pi/512
   cos[155]  =  6'b001001;     //155pi/512
   sin[156]  =  6'b110011;     //156pi/512
   cos[156]  =  6'b001001;     //156pi/512
   sin[157]  =  6'b110011;     //157pi/512
   cos[157]  =  6'b001001;     //157pi/512
   sin[158]  =  6'b110011;     //158pi/512
   cos[158]  =  6'b001001;     //158pi/512
   sin[159]  =  6'b110011;     //159pi/512
   cos[159]  =  6'b001000;     //159pi/512
   sin[160]  =  6'b110011;     //160pi/512
   cos[160]  =  6'b001000;     //160pi/512
   sin[161]  =  6'b110011;     //161pi/512
   cos[161]  =  6'b001000;     //161pi/512
   sin[162]  =  6'b110011;     //162pi/512
   cos[162]  =  6'b001000;     //162pi/512
   sin[163]  =  6'b110011;     //163pi/512
   cos[163]  =  6'b001000;     //163pi/512
   sin[164]  =  6'b110010;     //164pi/512
   cos[164]  =  6'b001000;     //164pi/512
   sin[165]  =  6'b110010;     //165pi/512
   cos[165]  =  6'b001000;     //165pi/512
   sin[166]  =  6'b110010;     //166pi/512
   cos[166]  =  6'b001000;     //166pi/512
   sin[167]  =  6'b110010;     //167pi/512
   cos[167]  =  6'b001000;     //167pi/512
   sin[168]  =  6'b110010;     //168pi/512
   cos[168]  =  6'b001000;     //168pi/512
   sin[169]  =  6'b110010;     //169pi/512
   cos[169]  =  6'b001000;     //169pi/512
   sin[170]  =  6'b110010;     //170pi/512
   cos[170]  =  6'b001000;     //170pi/512
   sin[171]  =  6'b110010;     //171pi/512
   cos[171]  =  6'b000111;     //171pi/512
   sin[172]  =  6'b110010;     //172pi/512
   cos[172]  =  6'b000111;     //172pi/512
   sin[173]  =  6'b110010;     //173pi/512
   cos[173]  =  6'b000111;     //173pi/512
   sin[174]  =  6'b110010;     //174pi/512
   cos[174]  =  6'b000111;     //174pi/512
   sin[175]  =  6'b110010;     //175pi/512
   cos[175]  =  6'b000111;     //175pi/512
   sin[176]  =  6'b110010;     //176pi/512
   cos[176]  =  6'b000111;     //176pi/512
   sin[177]  =  6'b110010;     //177pi/512
   cos[177]  =  6'b000111;     //177pi/512
   sin[178]  =  6'b110010;     //178pi/512
   cos[178]  =  6'b000111;     //178pi/512
   sin[179]  =  6'b110010;     //179pi/512
   cos[179]  =  6'b000111;     //179pi/512
   sin[180]  =  6'b110010;     //180pi/512
   cos[180]  =  6'b000111;     //180pi/512
   sin[181]  =  6'b110010;     //181pi/512
   cos[181]  =  6'b000111;     //181pi/512
   sin[182]  =  6'b110010;     //182pi/512
   cos[182]  =  6'b000111;     //182pi/512
   sin[183]  =  6'b110010;     //183pi/512
   cos[183]  =  6'b000110;     //183pi/512
   sin[184]  =  6'b110010;     //184pi/512
   cos[184]  =  6'b000110;     //184pi/512
   sin[185]  =  6'b110001;     //185pi/512
   cos[185]  =  6'b000110;     //185pi/512
   sin[186]  =  6'b110001;     //186pi/512
   cos[186]  =  6'b000110;     //186pi/512
   sin[187]  =  6'b110001;     //187pi/512
   cos[187]  =  6'b000110;     //187pi/512
   sin[188]  =  6'b110001;     //188pi/512
   cos[188]  =  6'b000110;     //188pi/512
   sin[189]  =  6'b110001;     //189pi/512
   cos[189]  =  6'b000110;     //189pi/512
   sin[190]  =  6'b110001;     //190pi/512
   cos[190]  =  6'b000110;     //190pi/512
   sin[191]  =  6'b110001;     //191pi/512
   cos[191]  =  6'b000110;     //191pi/512
   sin[192]  =  6'b110001;     //192pi/512
   cos[192]  =  6'b000110;     //192pi/512
   sin[193]  =  6'b110001;     //193pi/512
   cos[193]  =  6'b000110;     //193pi/512
   sin[194]  =  6'b110001;     //194pi/512
   cos[194]  =  6'b000101;     //194pi/512
   sin[195]  =  6'b110001;     //195pi/512
   cos[195]  =  6'b000101;     //195pi/512
   sin[196]  =  6'b110001;     //196pi/512
   cos[196]  =  6'b000101;     //196pi/512
   sin[197]  =  6'b110001;     //197pi/512
   cos[197]  =  6'b000101;     //197pi/512
   sin[198]  =  6'b110001;     //198pi/512
   cos[198]  =  6'b000101;     //198pi/512
   sin[199]  =  6'b110001;     //199pi/512
   cos[199]  =  6'b000101;     //199pi/512
   sin[200]  =  6'b110001;     //200pi/512
   cos[200]  =  6'b000101;     //200pi/512
   sin[201]  =  6'b110001;     //201pi/512
   cos[201]  =  6'b000101;     //201pi/512
   sin[202]  =  6'b110001;     //202pi/512
   cos[202]  =  6'b000101;     //202pi/512
   sin[203]  =  6'b110001;     //203pi/512
   cos[203]  =  6'b000101;     //203pi/512
   sin[204]  =  6'b110001;     //204pi/512
   cos[204]  =  6'b000101;     //204pi/512
   sin[205]  =  6'b110001;     //205pi/512
   cos[205]  =  6'b000100;     //205pi/512
   sin[206]  =  6'b110001;     //206pi/512
   cos[206]  =  6'b000100;     //206pi/512
   sin[207]  =  6'b110001;     //207pi/512
   cos[207]  =  6'b000100;     //207pi/512
   sin[208]  =  6'b110001;     //208pi/512
   cos[208]  =  6'b000100;     //208pi/512
   sin[209]  =  6'b110001;     //209pi/512
   cos[209]  =  6'b000100;     //209pi/512
   sin[210]  =  6'b110001;     //210pi/512
   cos[210]  =  6'b000100;     //210pi/512
   sin[211]  =  6'b110001;     //211pi/512
   cos[211]  =  6'b000100;     //211pi/512
   sin[212]  =  6'b110001;     //212pi/512
   cos[212]  =  6'b000100;     //212pi/512
   sin[213]  =  6'b110001;     //213pi/512
   cos[213]  =  6'b000100;     //213pi/512
   sin[214]  =  6'b110001;     //214pi/512
   cos[214]  =  6'b000100;     //214pi/512
   sin[215]  =  6'b110001;     //215pi/512
   cos[215]  =  6'b000011;     //215pi/512
   sin[216]  =  6'b110000;     //216pi/512
   cos[216]  =  6'b000011;     //216pi/512
   sin[217]  =  6'b110000;     //217pi/512
   cos[217]  =  6'b000011;     //217pi/512
   sin[218]  =  6'b110000;     //218pi/512
   cos[218]  =  6'b000011;     //218pi/512
   sin[219]  =  6'b110000;     //219pi/512
   cos[219]  =  6'b000011;     //219pi/512
   sin[220]  =  6'b110000;     //220pi/512
   cos[220]  =  6'b000011;     //220pi/512
   sin[221]  =  6'b110000;     //221pi/512
   cos[221]  =  6'b000011;     //221pi/512
   sin[222]  =  6'b110000;     //222pi/512
   cos[222]  =  6'b000011;     //222pi/512
   sin[223]  =  6'b110000;     //223pi/512
   cos[223]  =  6'b000011;     //223pi/512
   sin[224]  =  6'b110000;     //224pi/512
   cos[224]  =  6'b000011;     //224pi/512
   sin[225]  =  6'b110000;     //225pi/512
   cos[225]  =  6'b000011;     //225pi/512
   sin[226]  =  6'b110000;     //226pi/512
   cos[226]  =  6'b000010;     //226pi/512
   sin[227]  =  6'b110000;     //227pi/512
   cos[227]  =  6'b000010;     //227pi/512
   sin[228]  =  6'b110000;     //228pi/512
   cos[228]  =  6'b000010;     //228pi/512
   sin[229]  =  6'b110000;     //229pi/512
   cos[229]  =  6'b000010;     //229pi/512
   sin[230]  =  6'b110000;     //230pi/512
   cos[230]  =  6'b000010;     //230pi/512
   sin[231]  =  6'b110000;     //231pi/512
   cos[231]  =  6'b000010;     //231pi/512
   sin[232]  =  6'b110000;     //232pi/512
   cos[232]  =  6'b000010;     //232pi/512
   sin[233]  =  6'b110000;     //233pi/512
   cos[233]  =  6'b000010;     //233pi/512
   sin[234]  =  6'b110000;     //234pi/512
   cos[234]  =  6'b000010;     //234pi/512
   sin[235]  =  6'b110000;     //235pi/512
   cos[235]  =  6'b000010;     //235pi/512
   sin[236]  =  6'b110000;     //236pi/512
   cos[236]  =  6'b000001;     //236pi/512
   sin[237]  =  6'b110000;     //237pi/512
   cos[237]  =  6'b000001;     //237pi/512
   sin[238]  =  6'b110000;     //238pi/512
   cos[238]  =  6'b000001;     //238pi/512
   sin[239]  =  6'b110000;     //239pi/512
   cos[239]  =  6'b000001;     //239pi/512
   sin[240]  =  6'b110000;     //240pi/512
   cos[240]  =  6'b000001;     //240pi/512
   sin[241]  =  6'b110000;     //241pi/512
   cos[241]  =  6'b000001;     //241pi/512
   sin[242]  =  6'b110000;     //242pi/512
   cos[242]  =  6'b000001;     //242pi/512
   sin[243]  =  6'b110000;     //243pi/512
   cos[243]  =  6'b000001;     //243pi/512
   sin[244]  =  6'b110000;     //244pi/512
   cos[244]  =  6'b000001;     //244pi/512
   sin[245]  =  6'b110000;     //245pi/512
   cos[245]  =  6'b000001;     //245pi/512
   sin[246]  =  6'b110000;     //246pi/512
   cos[246]  =  6'b000000;     //246pi/512
   sin[247]  =  6'b110000;     //247pi/512
   cos[247]  =  6'b000000;     //247pi/512
   sin[248]  =  6'b110000;     //248pi/512
   cos[248]  =  6'b000000;     //248pi/512
   sin[249]  =  6'b110000;     //249pi/512
   cos[249]  =  6'b000000;     //249pi/512
   sin[250]  =  6'b110000;     //250pi/512
   cos[250]  =  6'b000000;     //250pi/512
   sin[251]  =  6'b110000;     //251pi/512
   cos[251]  =  6'b000000;     //251pi/512
   sin[252]  =  6'b110000;     //252pi/512
   cos[252]  =  6'b000000;     //252pi/512
   sin[253]  =  6'b110000;     //253pi/512
   cos[253]  =  6'b000000;     //253pi/512
   sin[254]  =  6'b110000;     //254pi/512
   cos[254]  =  6'b000000;     //254pi/512
   sin[255]  =  6'b110000;     //255pi/512
   cos[255]  =  6'b000000;     //255pi/512
   sin[256]  =  6'b110000;     //256pi/512
   cos[256]  =  6'b000000;     //256pi/512
   sin[257]  =  6'b110000;     //257pi/512
   cos[257]  =  6'b000000;     //257pi/512
   sin[258]  =  6'b110000;     //258pi/512
   cos[258]  =  6'b000000;     //258pi/512
   sin[259]  =  6'b110000;     //259pi/512
   cos[259]  =  6'b000000;     //259pi/512
   sin[260]  =  6'b110000;     //260pi/512
   cos[260]  =  6'b000000;     //260pi/512
   sin[261]  =  6'b110000;     //261pi/512
   cos[261]  =  6'b000000;     //261pi/512
   sin[262]  =  6'b110000;     //262pi/512
   cos[262]  =  6'b111111;     //262pi/512
   sin[263]  =  6'b110000;     //263pi/512
   cos[263]  =  6'b111111;     //263pi/512
   sin[264]  =  6'b110000;     //264pi/512
   cos[264]  =  6'b111111;     //264pi/512
   sin[265]  =  6'b110000;     //265pi/512
   cos[265]  =  6'b111111;     //265pi/512
   sin[266]  =  6'b110000;     //266pi/512
   cos[266]  =  6'b111111;     //266pi/512
   sin[267]  =  6'b110000;     //267pi/512
   cos[267]  =  6'b111111;     //267pi/512
   sin[268]  =  6'b110000;     //268pi/512
   cos[268]  =  6'b111111;     //268pi/512
   sin[269]  =  6'b110000;     //269pi/512
   cos[269]  =  6'b111111;     //269pi/512
   sin[270]  =  6'b110000;     //270pi/512
   cos[270]  =  6'b111111;     //270pi/512
   sin[271]  =  6'b110000;     //271pi/512
   cos[271]  =  6'b111111;     //271pi/512
   sin[272]  =  6'b110000;     //272pi/512
   cos[272]  =  6'b111110;     //272pi/512
   sin[273]  =  6'b110000;     //273pi/512
   cos[273]  =  6'b111110;     //273pi/512
   sin[274]  =  6'b110000;     //274pi/512
   cos[274]  =  6'b111110;     //274pi/512
   sin[275]  =  6'b110000;     //275pi/512
   cos[275]  =  6'b111110;     //275pi/512
   sin[276]  =  6'b110000;     //276pi/512
   cos[276]  =  6'b111110;     //276pi/512
   sin[277]  =  6'b110000;     //277pi/512
   cos[277]  =  6'b111110;     //277pi/512
   sin[278]  =  6'b110000;     //278pi/512
   cos[278]  =  6'b111110;     //278pi/512
   sin[279]  =  6'b110000;     //279pi/512
   cos[279]  =  6'b111110;     //279pi/512
   sin[280]  =  6'b110000;     //280pi/512
   cos[280]  =  6'b111110;     //280pi/512
   sin[281]  =  6'b110000;     //281pi/512
   cos[281]  =  6'b111110;     //281pi/512
   sin[282]  =  6'b110000;     //282pi/512
   cos[282]  =  6'b111101;     //282pi/512
   sin[283]  =  6'b110000;     //283pi/512
   cos[283]  =  6'b111101;     //283pi/512
   sin[284]  =  6'b110000;     //284pi/512
   cos[284]  =  6'b111101;     //284pi/512
   sin[285]  =  6'b110000;     //285pi/512
   cos[285]  =  6'b111101;     //285pi/512
   sin[286]  =  6'b110000;     //286pi/512
   cos[286]  =  6'b111101;     //286pi/512
   sin[287]  =  6'b110000;     //287pi/512
   cos[287]  =  6'b111101;     //287pi/512
   sin[288]  =  6'b110000;     //288pi/512
   cos[288]  =  6'b111101;     //288pi/512
   sin[289]  =  6'b110000;     //289pi/512
   cos[289]  =  6'b111101;     //289pi/512
   sin[290]  =  6'b110000;     //290pi/512
   cos[290]  =  6'b111101;     //290pi/512
   sin[291]  =  6'b110000;     //291pi/512
   cos[291]  =  6'b111101;     //291pi/512
   sin[292]  =  6'b110000;     //292pi/512
   cos[292]  =  6'b111100;     //292pi/512
   sin[293]  =  6'b110000;     //293pi/512
   cos[293]  =  6'b111100;     //293pi/512
   sin[294]  =  6'b110000;     //294pi/512
   cos[294]  =  6'b111100;     //294pi/512
   sin[295]  =  6'b110000;     //295pi/512
   cos[295]  =  6'b111100;     //295pi/512
   sin[296]  =  6'b110000;     //296pi/512
   cos[296]  =  6'b111100;     //296pi/512
   sin[297]  =  6'b110001;     //297pi/512
   cos[297]  =  6'b111100;     //297pi/512
   sin[298]  =  6'b110001;     //298pi/512
   cos[298]  =  6'b111100;     //298pi/512
   sin[299]  =  6'b110001;     //299pi/512
   cos[299]  =  6'b111100;     //299pi/512
   sin[300]  =  6'b110001;     //300pi/512
   cos[300]  =  6'b111100;     //300pi/512
   sin[301]  =  6'b110001;     //301pi/512
   cos[301]  =  6'b111100;     //301pi/512
   sin[302]  =  6'b110001;     //302pi/512
   cos[302]  =  6'b111100;     //302pi/512
   sin[303]  =  6'b110001;     //303pi/512
   cos[303]  =  6'b111011;     //303pi/512
   sin[304]  =  6'b110001;     //304pi/512
   cos[304]  =  6'b111011;     //304pi/512
   sin[305]  =  6'b110001;     //305pi/512
   cos[305]  =  6'b111011;     //305pi/512
   sin[306]  =  6'b110001;     //306pi/512
   cos[306]  =  6'b111011;     //306pi/512
   sin[307]  =  6'b110001;     //307pi/512
   cos[307]  =  6'b111011;     //307pi/512
   sin[308]  =  6'b110001;     //308pi/512
   cos[308]  =  6'b111011;     //308pi/512
   sin[309]  =  6'b110001;     //309pi/512
   cos[309]  =  6'b111011;     //309pi/512
   sin[310]  =  6'b110001;     //310pi/512
   cos[310]  =  6'b111011;     //310pi/512
   sin[311]  =  6'b110001;     //311pi/512
   cos[311]  =  6'b111011;     //311pi/512
   sin[312]  =  6'b110001;     //312pi/512
   cos[312]  =  6'b111011;     //312pi/512
   sin[313]  =  6'b110001;     //313pi/512
   cos[313]  =  6'b111011;     //313pi/512
   sin[314]  =  6'b110001;     //314pi/512
   cos[314]  =  6'b111010;     //314pi/512
   sin[315]  =  6'b110001;     //315pi/512
   cos[315]  =  6'b111010;     //315pi/512
   sin[316]  =  6'b110001;     //316pi/512
   cos[316]  =  6'b111010;     //316pi/512
   sin[317]  =  6'b110001;     //317pi/512
   cos[317]  =  6'b111010;     //317pi/512
   sin[318]  =  6'b110001;     //318pi/512
   cos[318]  =  6'b111010;     //318pi/512
   sin[319]  =  6'b110001;     //319pi/512
   cos[319]  =  6'b111010;     //319pi/512
   sin[320]  =  6'b110001;     //320pi/512
   cos[320]  =  6'b111010;     //320pi/512
   sin[321]  =  6'b110001;     //321pi/512
   cos[321]  =  6'b111010;     //321pi/512
   sin[322]  =  6'b110001;     //322pi/512
   cos[322]  =  6'b111010;     //322pi/512
   sin[323]  =  6'b110001;     //323pi/512
   cos[323]  =  6'b111010;     //323pi/512
   sin[324]  =  6'b110001;     //324pi/512
   cos[324]  =  6'b111010;     //324pi/512
   sin[325]  =  6'b110001;     //325pi/512
   cos[325]  =  6'b111001;     //325pi/512
   sin[326]  =  6'b110001;     //326pi/512
   cos[326]  =  6'b111001;     //326pi/512
   sin[327]  =  6'b110001;     //327pi/512
   cos[327]  =  6'b111001;     //327pi/512
   sin[328]  =  6'b110010;     //328pi/512
   cos[328]  =  6'b111001;     //328pi/512
   sin[329]  =  6'b110010;     //329pi/512
   cos[329]  =  6'b111001;     //329pi/512
   sin[330]  =  6'b110010;     //330pi/512
   cos[330]  =  6'b111001;     //330pi/512
   sin[331]  =  6'b110010;     //331pi/512
   cos[331]  =  6'b111001;     //331pi/512
   sin[332]  =  6'b110010;     //332pi/512
   cos[332]  =  6'b111001;     //332pi/512
   sin[333]  =  6'b110010;     //333pi/512
   cos[333]  =  6'b111001;     //333pi/512
   sin[334]  =  6'b110010;     //334pi/512
   cos[334]  =  6'b111001;     //334pi/512
   sin[335]  =  6'b110010;     //335pi/512
   cos[335]  =  6'b111001;     //335pi/512
   sin[336]  =  6'b110010;     //336pi/512
   cos[336]  =  6'b111000;     //336pi/512
   sin[337]  =  6'b110010;     //337pi/512
   cos[337]  =  6'b111000;     //337pi/512
   sin[338]  =  6'b110010;     //338pi/512
   cos[338]  =  6'b111000;     //338pi/512
   sin[339]  =  6'b110010;     //339pi/512
   cos[339]  =  6'b111000;     //339pi/512
   sin[340]  =  6'b110010;     //340pi/512
   cos[340]  =  6'b111000;     //340pi/512
   sin[341]  =  6'b110010;     //341pi/512
   cos[341]  =  6'b111000;     //341pi/512
   sin[342]  =  6'b110010;     //342pi/512
   cos[342]  =  6'b111000;     //342pi/512
   sin[343]  =  6'b110010;     //343pi/512
   cos[343]  =  6'b111000;     //343pi/512
   sin[344]  =  6'b110010;     //344pi/512
   cos[344]  =  6'b111000;     //344pi/512
   sin[345]  =  6'b110010;     //345pi/512
   cos[345]  =  6'b111000;     //345pi/512
   sin[346]  =  6'b110010;     //346pi/512
   cos[346]  =  6'b111000;     //346pi/512
   sin[347]  =  6'b110010;     //347pi/512
   cos[347]  =  6'b111000;     //347pi/512
   sin[348]  =  6'b110010;     //348pi/512
   cos[348]  =  6'b110111;     //348pi/512
   sin[349]  =  6'b110011;     //349pi/512
   cos[349]  =  6'b110111;     //349pi/512
   sin[350]  =  6'b110011;     //350pi/512
   cos[350]  =  6'b110111;     //350pi/512
   sin[351]  =  6'b110011;     //351pi/512
   cos[351]  =  6'b110111;     //351pi/512
   sin[352]  =  6'b110011;     //352pi/512
   cos[352]  =  6'b110111;     //352pi/512
   sin[353]  =  6'b110011;     //353pi/512
   cos[353]  =  6'b110111;     //353pi/512
   sin[354]  =  6'b110011;     //354pi/512
   cos[354]  =  6'b110111;     //354pi/512
   sin[355]  =  6'b110011;     //355pi/512
   cos[355]  =  6'b110111;     //355pi/512
   sin[356]  =  6'b110011;     //356pi/512
   cos[356]  =  6'b110111;     //356pi/512
   sin[357]  =  6'b110011;     //357pi/512
   cos[357]  =  6'b110111;     //357pi/512
   sin[358]  =  6'b110011;     //358pi/512
   cos[358]  =  6'b110111;     //358pi/512
   sin[359]  =  6'b110011;     //359pi/512
   cos[359]  =  6'b110111;     //359pi/512
   sin[360]  =  6'b110011;     //360pi/512
   cos[360]  =  6'b110110;     //360pi/512
   sin[361]  =  6'b110011;     //361pi/512
   cos[361]  =  6'b110110;     //361pi/512
   sin[362]  =  6'b110011;     //362pi/512
   cos[362]  =  6'b110110;     //362pi/512
   sin[363]  =  6'b110011;     //363pi/512
   cos[363]  =  6'b110110;     //363pi/512
   sin[364]  =  6'b110011;     //364pi/512
   cos[364]  =  6'b110110;     //364pi/512
   sin[365]  =  6'b110011;     //365pi/512
   cos[365]  =  6'b110110;     //365pi/512
   sin[366]  =  6'b110100;     //366pi/512
   cos[366]  =  6'b110110;     //366pi/512
   sin[367]  =  6'b110100;     //367pi/512
   cos[367]  =  6'b110110;     //367pi/512
   sin[368]  =  6'b110100;     //368pi/512
   cos[368]  =  6'b110110;     //368pi/512
   sin[369]  =  6'b110100;     //369pi/512
   cos[369]  =  6'b110110;     //369pi/512
   sin[370]  =  6'b110100;     //370pi/512
   cos[370]  =  6'b110110;     //370pi/512
   sin[371]  =  6'b110100;     //371pi/512
   cos[371]  =  6'b110110;     //371pi/512
   sin[372]  =  6'b110100;     //372pi/512
   cos[372]  =  6'b110110;     //372pi/512
   sin[373]  =  6'b110100;     //373pi/512
   cos[373]  =  6'b110101;     //373pi/512
   sin[374]  =  6'b110100;     //374pi/512
   cos[374]  =  6'b110101;     //374pi/512
   sin[375]  =  6'b110100;     //375pi/512
   cos[375]  =  6'b110101;     //375pi/512
   sin[376]  =  6'b110100;     //376pi/512
   cos[376]  =  6'b110101;     //376pi/512
   sin[377]  =  6'b110100;     //377pi/512
   cos[377]  =  6'b110101;     //377pi/512
   sin[378]  =  6'b110100;     //378pi/512
   cos[378]  =  6'b110101;     //378pi/512
   sin[379]  =  6'b110100;     //379pi/512
   cos[379]  =  6'b110101;     //379pi/512
   sin[380]  =  6'b110100;     //380pi/512
   cos[380]  =  6'b110101;     //380pi/512
   sin[381]  =  6'b110100;     //381pi/512
   cos[381]  =  6'b110101;     //381pi/512
   sin[382]  =  6'b110101;     //382pi/512
   cos[382]  =  6'b110101;     //382pi/512
   sin[383]  =  6'b110101;     //383pi/512
   cos[383]  =  6'b110101;     //383pi/512
   sin[384]  =  6'b110101;     //384pi/512
   cos[384]  =  6'b110101;     //384pi/512
   sin[385]  =  6'b110101;     //385pi/512
   cos[385]  =  6'b110101;     //385pi/512
   sin[386]  =  6'b110101;     //386pi/512
   cos[386]  =  6'b110101;     //386pi/512
   sin[387]  =  6'b110101;     //387pi/512
   cos[387]  =  6'b110100;     //387pi/512
   sin[388]  =  6'b110101;     //388pi/512
   cos[388]  =  6'b110100;     //388pi/512
   sin[389]  =  6'b110101;     //389pi/512
   cos[389]  =  6'b110100;     //389pi/512
   sin[390]  =  6'b110101;     //390pi/512
   cos[390]  =  6'b110100;     //390pi/512
   sin[391]  =  6'b110101;     //391pi/512
   cos[391]  =  6'b110100;     //391pi/512
   sin[392]  =  6'b110101;     //392pi/512
   cos[392]  =  6'b110100;     //392pi/512
   sin[393]  =  6'b110101;     //393pi/512
   cos[393]  =  6'b110100;     //393pi/512
   sin[394]  =  6'b110101;     //394pi/512
   cos[394]  =  6'b110100;     //394pi/512
   sin[395]  =  6'b110101;     //395pi/512
   cos[395]  =  6'b110100;     //395pi/512
   sin[396]  =  6'b110110;     //396pi/512
   cos[396]  =  6'b110100;     //396pi/512
   sin[397]  =  6'b110110;     //397pi/512
   cos[397]  =  6'b110100;     //397pi/512
   sin[398]  =  6'b110110;     //398pi/512
   cos[398]  =  6'b110100;     //398pi/512
   sin[399]  =  6'b110110;     //399pi/512
   cos[399]  =  6'b110100;     //399pi/512
   sin[400]  =  6'b110110;     //400pi/512
   cos[400]  =  6'b110100;     //400pi/512
   sin[401]  =  6'b110110;     //401pi/512
   cos[401]  =  6'b110100;     //401pi/512
   sin[402]  =  6'b110110;     //402pi/512
   cos[402]  =  6'b110100;     //402pi/512
   sin[403]  =  6'b110110;     //403pi/512
   cos[403]  =  6'b110011;     //403pi/512
   sin[404]  =  6'b110110;     //404pi/512
   cos[404]  =  6'b110011;     //404pi/512
   sin[405]  =  6'b110110;     //405pi/512
   cos[405]  =  6'b110011;     //405pi/512
   sin[406]  =  6'b110110;     //406pi/512
   cos[406]  =  6'b110011;     //406pi/512
   sin[407]  =  6'b110110;     //407pi/512
   cos[407]  =  6'b110011;     //407pi/512
   sin[408]  =  6'b110110;     //408pi/512
   cos[408]  =  6'b110011;     //408pi/512
   sin[409]  =  6'b110111;     //409pi/512
   cos[409]  =  6'b110011;     //409pi/512
   sin[410]  =  6'b110111;     //410pi/512
   cos[410]  =  6'b110011;     //410pi/512
   sin[411]  =  6'b110111;     //411pi/512
   cos[411]  =  6'b110011;     //411pi/512
   sin[412]  =  6'b110111;     //412pi/512
   cos[412]  =  6'b110011;     //412pi/512
   sin[413]  =  6'b110111;     //413pi/512
   cos[413]  =  6'b110011;     //413pi/512
   sin[414]  =  6'b110111;     //414pi/512
   cos[414]  =  6'b110011;     //414pi/512
   sin[415]  =  6'b110111;     //415pi/512
   cos[415]  =  6'b110011;     //415pi/512
   sin[416]  =  6'b110111;     //416pi/512
   cos[416]  =  6'b110011;     //416pi/512
   sin[417]  =  6'b110111;     //417pi/512
   cos[417]  =  6'b110011;     //417pi/512
   sin[418]  =  6'b110111;     //418pi/512
   cos[418]  =  6'b110011;     //418pi/512
   sin[419]  =  6'b110111;     //419pi/512
   cos[419]  =  6'b110011;     //419pi/512
   sin[420]  =  6'b110111;     //420pi/512
   cos[420]  =  6'b110010;     //420pi/512
   sin[421]  =  6'b111000;     //421pi/512
   cos[421]  =  6'b110010;     //421pi/512
   sin[422]  =  6'b111000;     //422pi/512
   cos[422]  =  6'b110010;     //422pi/512
   sin[423]  =  6'b111000;     //423pi/512
   cos[423]  =  6'b110010;     //423pi/512
   sin[424]  =  6'b111000;     //424pi/512
   cos[424]  =  6'b110010;     //424pi/512
   sin[425]  =  6'b111000;     //425pi/512
   cos[425]  =  6'b110010;     //425pi/512
   sin[426]  =  6'b111000;     //426pi/512
   cos[426]  =  6'b110010;     //426pi/512
   sin[427]  =  6'b111000;     //427pi/512
   cos[427]  =  6'b110010;     //427pi/512
   sin[428]  =  6'b111000;     //428pi/512
   cos[428]  =  6'b110010;     //428pi/512
   sin[429]  =  6'b111000;     //429pi/512
   cos[429]  =  6'b110010;     //429pi/512
   sin[430]  =  6'b111000;     //430pi/512
   cos[430]  =  6'b110010;     //430pi/512
   sin[431]  =  6'b111000;     //431pi/512
   cos[431]  =  6'b110010;     //431pi/512
   sin[432]  =  6'b111000;     //432pi/512
   cos[432]  =  6'b110010;     //432pi/512
   sin[433]  =  6'b111001;     //433pi/512
   cos[433]  =  6'b110010;     //433pi/512
   sin[434]  =  6'b111001;     //434pi/512
   cos[434]  =  6'b110010;     //434pi/512
   sin[435]  =  6'b111001;     //435pi/512
   cos[435]  =  6'b110010;     //435pi/512
   sin[436]  =  6'b111001;     //436pi/512
   cos[436]  =  6'b110010;     //436pi/512
   sin[437]  =  6'b111001;     //437pi/512
   cos[437]  =  6'b110010;     //437pi/512
   sin[438]  =  6'b111001;     //438pi/512
   cos[438]  =  6'b110010;     //438pi/512
   sin[439]  =  6'b111001;     //439pi/512
   cos[439]  =  6'b110010;     //439pi/512
   sin[440]  =  6'b111001;     //440pi/512
   cos[440]  =  6'b110010;     //440pi/512
   sin[441]  =  6'b111001;     //441pi/512
   cos[441]  =  6'b110001;     //441pi/512
   sin[442]  =  6'b111001;     //442pi/512
   cos[442]  =  6'b110001;     //442pi/512
   sin[443]  =  6'b111001;     //443pi/512
   cos[443]  =  6'b110001;     //443pi/512
   sin[444]  =  6'b111010;     //444pi/512
   cos[444]  =  6'b110001;     //444pi/512
   sin[445]  =  6'b111010;     //445pi/512
   cos[445]  =  6'b110001;     //445pi/512
   sin[446]  =  6'b111010;     //446pi/512
   cos[446]  =  6'b110001;     //446pi/512
   sin[447]  =  6'b111010;     //447pi/512
   cos[447]  =  6'b110001;     //447pi/512
   sin[448]  =  6'b111010;     //448pi/512
   cos[448]  =  6'b110001;     //448pi/512
   sin[449]  =  6'b111010;     //449pi/512
   cos[449]  =  6'b110001;     //449pi/512
   sin[450]  =  6'b111010;     //450pi/512
   cos[450]  =  6'b110001;     //450pi/512
   sin[451]  =  6'b111010;     //451pi/512
   cos[451]  =  6'b110001;     //451pi/512
   sin[452]  =  6'b111010;     //452pi/512
   cos[452]  =  6'b110001;     //452pi/512
   sin[453]  =  6'b111010;     //453pi/512
   cos[453]  =  6'b110001;     //453pi/512
   sin[454]  =  6'b111010;     //454pi/512
   cos[454]  =  6'b110001;     //454pi/512
   sin[455]  =  6'b111011;     //455pi/512
   cos[455]  =  6'b110001;     //455pi/512
   sin[456]  =  6'b111011;     //456pi/512
   cos[456]  =  6'b110001;     //456pi/512
   sin[457]  =  6'b111011;     //457pi/512
   cos[457]  =  6'b110001;     //457pi/512
   sin[458]  =  6'b111011;     //458pi/512
   cos[458]  =  6'b110001;     //458pi/512
   sin[459]  =  6'b111011;     //459pi/512
   cos[459]  =  6'b110001;     //459pi/512
   sin[460]  =  6'b111011;     //460pi/512
   cos[460]  =  6'b110001;     //460pi/512
   sin[461]  =  6'b111011;     //461pi/512
   cos[461]  =  6'b110001;     //461pi/512
   sin[462]  =  6'b111011;     //462pi/512
   cos[462]  =  6'b110001;     //462pi/512
   sin[463]  =  6'b111011;     //463pi/512
   cos[463]  =  6'b110001;     //463pi/512
   sin[464]  =  6'b111011;     //464pi/512
   cos[464]  =  6'b110001;     //464pi/512
   sin[465]  =  6'b111011;     //465pi/512
   cos[465]  =  6'b110001;     //465pi/512
   sin[466]  =  6'b111100;     //466pi/512
   cos[466]  =  6'b110001;     //466pi/512
   sin[467]  =  6'b111100;     //467pi/512
   cos[467]  =  6'b110001;     //467pi/512
   sin[468]  =  6'b111100;     //468pi/512
   cos[468]  =  6'b110001;     //468pi/512
   sin[469]  =  6'b111100;     //469pi/512
   cos[469]  =  6'b110001;     //469pi/512
   sin[470]  =  6'b111100;     //470pi/512
   cos[470]  =  6'b110001;     //470pi/512
   sin[471]  =  6'b111100;     //471pi/512
   cos[471]  =  6'b110001;     //471pi/512
   sin[472]  =  6'b111100;     //472pi/512
   cos[472]  =  6'b110000;     //472pi/512
   sin[473]  =  6'b111100;     //473pi/512
   cos[473]  =  6'b110000;     //473pi/512
   sin[474]  =  6'b111100;     //474pi/512
   cos[474]  =  6'b110000;     //474pi/512
   sin[475]  =  6'b111100;     //475pi/512
   cos[475]  =  6'b110000;     //475pi/512
   sin[476]  =  6'b111100;     //476pi/512
   cos[476]  =  6'b110000;     //476pi/512
   sin[477]  =  6'b111101;     //477pi/512
   cos[477]  =  6'b110000;     //477pi/512
   sin[478]  =  6'b111101;     //478pi/512
   cos[478]  =  6'b110000;     //478pi/512
   sin[479]  =  6'b111101;     //479pi/512
   cos[479]  =  6'b110000;     //479pi/512
   sin[480]  =  6'b111101;     //480pi/512
   cos[480]  =  6'b110000;     //480pi/512
   sin[481]  =  6'b111101;     //481pi/512
   cos[481]  =  6'b110000;     //481pi/512
   sin[482]  =  6'b111101;     //482pi/512
   cos[482]  =  6'b110000;     //482pi/512
   sin[483]  =  6'b111101;     //483pi/512
   cos[483]  =  6'b110000;     //483pi/512
   sin[484]  =  6'b111101;     //484pi/512
   cos[484]  =  6'b110000;     //484pi/512
   sin[485]  =  6'b111101;     //485pi/512
   cos[485]  =  6'b110000;     //485pi/512
   sin[486]  =  6'b111101;     //486pi/512
   cos[486]  =  6'b110000;     //486pi/512
   sin[487]  =  6'b111110;     //487pi/512
   cos[487]  =  6'b110000;     //487pi/512
   sin[488]  =  6'b111110;     //488pi/512
   cos[488]  =  6'b110000;     //488pi/512
   sin[489]  =  6'b111110;     //489pi/512
   cos[489]  =  6'b110000;     //489pi/512
   sin[490]  =  6'b111110;     //490pi/512
   cos[490]  =  6'b110000;     //490pi/512
   sin[491]  =  6'b111110;     //491pi/512
   cos[491]  =  6'b110000;     //491pi/512
   sin[492]  =  6'b111110;     //492pi/512
   cos[492]  =  6'b110000;     //492pi/512
   sin[493]  =  6'b111110;     //493pi/512
   cos[493]  =  6'b110000;     //493pi/512
   sin[494]  =  6'b111110;     //494pi/512
   cos[494]  =  6'b110000;     //494pi/512
   sin[495]  =  6'b111110;     //495pi/512
   cos[495]  =  6'b110000;     //495pi/512
   sin[496]  =  6'b111110;     //496pi/512
   cos[496]  =  6'b110000;     //496pi/512
   sin[497]  =  6'b111111;     //497pi/512
   cos[497]  =  6'b110000;     //497pi/512
   sin[498]  =  6'b111111;     //498pi/512
   cos[498]  =  6'b110000;     //498pi/512
   sin[499]  =  6'b111111;     //499pi/512
   cos[499]  =  6'b110000;     //499pi/512
   sin[500]  =  6'b111111;     //500pi/512
   cos[500]  =  6'b110000;     //500pi/512
   sin[501]  =  6'b111111;     //501pi/512
   cos[501]  =  6'b110000;     //501pi/512
   sin[502]  =  6'b111111;     //502pi/512
   cos[502]  =  6'b110000;     //502pi/512
   sin[503]  =  6'b111111;     //503pi/512
   cos[503]  =  6'b110000;     //503pi/512
   sin[504]  =  6'b111111;     //504pi/512
   cos[504]  =  6'b110000;     //504pi/512
   sin[505]  =  6'b111111;     //505pi/512
   cos[505]  =  6'b110000;     //505pi/512
   sin[506]  =  6'b111111;     //506pi/512
   cos[506]  =  6'b110000;     //506pi/512
   sin[507]  =  6'b000000;     //507pi/512
   cos[507]  =  6'b110000;     //507pi/512
   sin[508]  =  6'b000000;     //508pi/512
   cos[508]  =  6'b110000;     //508pi/512
   sin[509]  =  6'b000000;     //509pi/512
   cos[509]  =  6'b110000;     //509pi/512
   sin[510]  =  6'b000000;     //510pi/512
   cos[510]  =  6'b110000;     //510pi/512
   sin[511]  =  6'b000000;     //511pi/512
   cos[511]  =  6'b110000;     //511pi/512
/////////////////////////////////////////////////////////
   m_sin[0]  =  6'b000000;     //0pi/512
   m_cos[0]  =  6'b010000;     //0pi/512
   m_sin[1]  =  6'b000000;     //1pi/512
   m_cos[1]  =  6'b001111;     //1pi/512
   m_sin[2]  =  6'b000000;     //2pi/512
   m_cos[2]  =  6'b001111;     //2pi/512
   m_sin[3]  =  6'b000000;     //3pi/512
   m_cos[3]  =  6'b001111;     //3pi/512
   m_sin[4]  =  6'b000000;     //4pi/512
   m_cos[4]  =  6'b001111;     //4pi/512
   m_sin[5]  =  6'b000000;     //5pi/512
   m_cos[5]  =  6'b001111;     //5pi/512
   m_sin[6]  =  6'b000000;     //6pi/512
   m_cos[6]  =  6'b001111;     //6pi/512
   m_sin[7]  =  6'b111111;     //7pi/512
   m_cos[7]  =  6'b001111;     //7pi/512
   m_sin[8]  =  6'b111111;     //8pi/512
   m_cos[8]  =  6'b001111;     //8pi/512
   m_sin[9]  =  6'b111111;     //9pi/512
   m_cos[9]  =  6'b001111;     //9pi/512
   m_sin[10]  =  6'b111111;     //10pi/512
   m_cos[10]  =  6'b001111;     //10pi/512
   m_sin[11]  =  6'b111111;     //11pi/512
   m_cos[11]  =  6'b001111;     //11pi/512
   m_sin[12]  =  6'b111111;     //12pi/512
   m_cos[12]  =  6'b001111;     //12pi/512
   m_sin[13]  =  6'b111111;     //13pi/512
   m_cos[13]  =  6'b001111;     //13pi/512
   m_sin[14]  =  6'b111111;     //14pi/512
   m_cos[14]  =  6'b001111;     //14pi/512
   m_sin[15]  =  6'b111111;     //15pi/512
   m_cos[15]  =  6'b001111;     //15pi/512
   m_sin[16]  =  6'b111111;     //16pi/512
   m_cos[16]  =  6'b001111;     //16pi/512
   m_sin[17]  =  6'b111111;     //17pi/512
   m_cos[17]  =  6'b001111;     //17pi/512
   m_sin[18]  =  6'b111111;     //18pi/512
   m_cos[18]  =  6'b001111;     //18pi/512
   m_sin[19]  =  6'b111111;     //19pi/512
   m_cos[19]  =  6'b001111;     //19pi/512
   m_sin[20]  =  6'b111110;     //20pi/512
   m_cos[20]  =  6'b001111;     //20pi/512
   m_sin[21]  =  6'b111110;     //21pi/512
   m_cos[21]  =  6'b001111;     //21pi/512
   m_sin[22]  =  6'b111110;     //22pi/512
   m_cos[22]  =  6'b001111;     //22pi/512
   m_sin[23]  =  6'b111110;     //23pi/512
   m_cos[23]  =  6'b001111;     //23pi/512
   m_sin[24]  =  6'b111110;     //24pi/512
   m_cos[24]  =  6'b001111;     //24pi/512
   m_sin[25]  =  6'b111110;     //25pi/512
   m_cos[25]  =  6'b001111;     //25pi/512
   m_sin[26]  =  6'b111110;     //26pi/512
   m_cos[26]  =  6'b001111;     //26pi/512
   m_sin[27]  =  6'b111110;     //27pi/512
   m_cos[27]  =  6'b001111;     //27pi/512
   m_sin[28]  =  6'b111110;     //28pi/512
   m_cos[28]  =  6'b001111;     //28pi/512
   m_sin[29]  =  6'b111110;     //29pi/512
   m_cos[29]  =  6'b001111;     //29pi/512
   m_sin[30]  =  6'b111110;     //30pi/512
   m_cos[30]  =  6'b001111;     //30pi/512
   m_sin[31]  =  6'b111110;     //31pi/512
   m_cos[31]  =  6'b001111;     //31pi/512
   m_sin[32]  =  6'b111101;     //32pi/512
   m_cos[32]  =  6'b001111;     //32pi/512
   m_sin[33]  =  6'b111101;     //33pi/512
   m_cos[33]  =  6'b001111;     //33pi/512
   m_sin[34]  =  6'b111101;     //34pi/512
   m_cos[34]  =  6'b001111;     //34pi/512
   m_sin[35]  =  6'b111101;     //35pi/512
   m_cos[35]  =  6'b001111;     //35pi/512
   m_sin[36]  =  6'b111101;     //36pi/512
   m_cos[36]  =  6'b001111;     //36pi/512
   m_sin[37]  =  6'b111101;     //37pi/512
   m_cos[37]  =  6'b001111;     //37pi/512
   m_sin[38]  =  6'b111101;     //38pi/512
   m_cos[38]  =  6'b001111;     //38pi/512
   m_sin[39]  =  6'b111101;     //39pi/512
   m_cos[39]  =  6'b001111;     //39pi/512
   m_sin[40]  =  6'b111101;     //40pi/512
   m_cos[40]  =  6'b001111;     //40pi/512
   m_sin[41]  =  6'b111101;     //41pi/512
   m_cos[41]  =  6'b001111;     //41pi/512
   m_sin[42]  =  6'b111101;     //42pi/512
   m_cos[42]  =  6'b001111;     //42pi/512
   m_sin[43]  =  6'b111101;     //43pi/512
   m_cos[43]  =  6'b001111;     //43pi/512
   m_sin[44]  =  6'b111101;     //44pi/512
   m_cos[44]  =  6'b001111;     //44pi/512
   m_sin[45]  =  6'b111100;     //45pi/512
   m_cos[45]  =  6'b001111;     //45pi/512
   m_sin[46]  =  6'b111100;     //46pi/512
   m_cos[46]  =  6'b001111;     //46pi/512
   m_sin[47]  =  6'b111100;     //47pi/512
   m_cos[47]  =  6'b001111;     //47pi/512
   m_sin[48]  =  6'b111100;     //48pi/512
   m_cos[48]  =  6'b001111;     //48pi/512
   m_sin[49]  =  6'b111100;     //49pi/512
   m_cos[49]  =  6'b001111;     //49pi/512
   m_sin[50]  =  6'b111100;     //50pi/512
   m_cos[50]  =  6'b001111;     //50pi/512
   m_sin[51]  =  6'b111100;     //51pi/512
   m_cos[51]  =  6'b001111;     //51pi/512
   m_sin[52]  =  6'b111100;     //52pi/512
   m_cos[52]  =  6'b001111;     //52pi/512
   m_sin[53]  =  6'b111100;     //53pi/512
   m_cos[53]  =  6'b001111;     //53pi/512
   m_sin[54]  =  6'b111100;     //54pi/512
   m_cos[54]  =  6'b001111;     //54pi/512
   m_sin[55]  =  6'b111100;     //55pi/512
   m_cos[55]  =  6'b001111;     //55pi/512
   m_sin[56]  =  6'b111100;     //56pi/512
   m_cos[56]  =  6'b001111;     //56pi/512
   m_sin[57]  =  6'b111100;     //57pi/512
   m_cos[57]  =  6'b001111;     //57pi/512
   m_sin[58]  =  6'b111100;     //58pi/512
   m_cos[58]  =  6'b001111;     //58pi/512
   m_sin[59]  =  6'b111011;     //59pi/512
   m_cos[59]  =  6'b001111;     //59pi/512
   m_sin[60]  =  6'b111011;     //60pi/512
   m_cos[60]  =  6'b001111;     //60pi/512
   m_sin[61]  =  6'b111011;     //61pi/512
   m_cos[61]  =  6'b001111;     //61pi/512
   m_sin[62]  =  6'b111011;     //62pi/512
   m_cos[62]  =  6'b001111;     //62pi/512
   m_sin[63]  =  6'b111011;     //63pi/512
   m_cos[63]  =  6'b001111;     //63pi/512
   m_sin[64]  =  6'b111011;     //64pi/512
   m_cos[64]  =  6'b001111;     //64pi/512
   m_sin[65]  =  6'b111011;     //65pi/512
   m_cos[65]  =  6'b001111;     //65pi/512
   m_sin[66]  =  6'b111011;     //66pi/512
   m_cos[66]  =  6'b001111;     //66pi/512
   m_sin[67]  =  6'b111011;     //67pi/512
   m_cos[67]  =  6'b001111;     //67pi/512
   m_sin[68]  =  6'b111011;     //68pi/512
   m_cos[68]  =  6'b001111;     //68pi/512
   m_sin[69]  =  6'b111011;     //69pi/512
   m_cos[69]  =  6'b001111;     //69pi/512
   m_sin[70]  =  6'b111011;     //70pi/512
   m_cos[70]  =  6'b001111;     //70pi/512
   m_sin[71]  =  6'b111011;     //71pi/512
   m_cos[71]  =  6'b001111;     //71pi/512
   m_sin[72]  =  6'b111010;     //72pi/512
   m_cos[72]  =  6'b001111;     //72pi/512
   m_sin[73]  =  6'b111010;     //73pi/512
   m_cos[73]  =  6'b001110;     //73pi/512
   m_sin[74]  =  6'b111010;     //74pi/512
   m_cos[74]  =  6'b001110;     //74pi/512
   m_sin[75]  =  6'b111010;     //75pi/512
   m_cos[75]  =  6'b001110;     //75pi/512
   m_sin[76]  =  6'b111010;     //76pi/512
   m_cos[76]  =  6'b001110;     //76pi/512
   m_sin[77]  =  6'b111010;     //77pi/512
   m_cos[77]  =  6'b001110;     //77pi/512
   m_sin[78]  =  6'b111010;     //78pi/512
   m_cos[78]  =  6'b001110;     //78pi/512
   m_sin[79]  =  6'b111010;     //79pi/512
   m_cos[79]  =  6'b001110;     //79pi/512
   m_sin[80]  =  6'b111010;     //80pi/512
   m_cos[80]  =  6'b001110;     //80pi/512
   m_sin[81]  =  6'b111010;     //81pi/512
   m_cos[81]  =  6'b001110;     //81pi/512
   m_sin[82]  =  6'b111010;     //82pi/512
   m_cos[82]  =  6'b001110;     //82pi/512
   m_sin[83]  =  6'b111010;     //83pi/512
   m_cos[83]  =  6'b001110;     //83pi/512
   m_sin[84]  =  6'b111010;     //84pi/512
   m_cos[84]  =  6'b001110;     //84pi/512
   m_sin[85]  =  6'b111010;     //85pi/512
   m_cos[85]  =  6'b001110;     //85pi/512
   m_sin[86]  =  6'b111001;     //86pi/512
   m_cos[86]  =  6'b001110;     //86pi/512
   m_sin[87]  =  6'b111001;     //87pi/512
   m_cos[87]  =  6'b001110;     //87pi/512
   m_sin[88]  =  6'b111001;     //88pi/512
   m_cos[88]  =  6'b001110;     //88pi/512
   m_sin[89]  =  6'b111001;     //89pi/512
   m_cos[89]  =  6'b001110;     //89pi/512
   m_sin[90]  =  6'b111001;     //90pi/512
   m_cos[90]  =  6'b001110;     //90pi/512
   m_sin[91]  =  6'b111001;     //91pi/512
   m_cos[91]  =  6'b001110;     //91pi/512
   m_sin[92]  =  6'b111001;     //92pi/512
   m_cos[92]  =  6'b001110;     //92pi/512
   m_sin[93]  =  6'b111001;     //93pi/512
   m_cos[93]  =  6'b001110;     //93pi/512
   m_sin[94]  =  6'b111001;     //94pi/512
   m_cos[94]  =  6'b001110;     //94pi/512
   m_sin[95]  =  6'b111001;     //95pi/512
   m_cos[95]  =  6'b001110;     //95pi/512
   m_sin[96]  =  6'b111001;     //96pi/512
   m_cos[96]  =  6'b001110;     //96pi/512
   m_sin[97]  =  6'b111001;     //97pi/512
   m_cos[97]  =  6'b001110;     //97pi/512
   m_sin[98]  =  6'b111001;     //98pi/512
   m_cos[98]  =  6'b001110;     //98pi/512
   m_sin[99]  =  6'b111001;     //99pi/512
   m_cos[99]  =  6'b001110;     //99pi/512
   m_sin[100]  =  6'b111000;     //100pi/512
   m_cos[100]  =  6'b001110;     //100pi/512
   m_sin[101]  =  6'b111000;     //101pi/512
   m_cos[101]  =  6'b001110;     //101pi/512
   m_sin[102]  =  6'b111000;     //102pi/512
   m_cos[102]  =  6'b001110;     //102pi/512
   m_sin[103]  =  6'b111000;     //103pi/512
   m_cos[103]  =  6'b001101;     //103pi/512
   m_sin[104]  =  6'b111000;     //104pi/512
   m_cos[104]  =  6'b001101;     //104pi/512
   m_sin[105]  =  6'b111000;     //105pi/512
   m_cos[105]  =  6'b001101;     //105pi/512
   m_sin[106]  =  6'b111000;     //106pi/512
   m_cos[106]  =  6'b001101;     //106pi/512
   m_sin[107]  =  6'b111000;     //107pi/512
   m_cos[107]  =  6'b001101;     //107pi/512
   m_sin[108]  =  6'b111000;     //108pi/512
   m_cos[108]  =  6'b001101;     //108pi/512
   m_sin[109]  =  6'b111000;     //109pi/512
   m_cos[109]  =  6'b001101;     //109pi/512
   m_sin[110]  =  6'b111000;     //110pi/512
   m_cos[110]  =  6'b001101;     //110pi/512
   m_sin[111]  =  6'b111000;     //111pi/512
   m_cos[111]  =  6'b001101;     //111pi/512
   m_sin[112]  =  6'b111000;     //112pi/512
   m_cos[112]  =  6'b001101;     //112pi/512
   m_sin[113]  =  6'b111000;     //113pi/512
   m_cos[113]  =  6'b001101;     //113pi/512
   m_sin[114]  =  6'b111000;     //114pi/512
   m_cos[114]  =  6'b001101;     //114pi/512
   m_sin[115]  =  6'b110111;     //115pi/512
   m_cos[115]  =  6'b001101;     //115pi/512
   m_sin[116]  =  6'b110111;     //116pi/512
   m_cos[116]  =  6'b001101;     //116pi/512
   m_sin[117]  =  6'b110111;     //117pi/512
   m_cos[117]  =  6'b001101;     //117pi/512
   m_sin[118]  =  6'b110111;     //118pi/512
   m_cos[118]  =  6'b001101;     //118pi/512
   m_sin[119]  =  6'b110111;     //119pi/512
   m_cos[119]  =  6'b001101;     //119pi/512
   m_sin[120]  =  6'b110111;     //120pi/512
   m_cos[120]  =  6'b001101;     //120pi/512
   m_sin[121]  =  6'b110111;     //121pi/512
   m_cos[121]  =  6'b001101;     //121pi/512
   m_sin[122]  =  6'b110111;     //122pi/512
   m_cos[122]  =  6'b001101;     //122pi/512
   m_sin[123]  =  6'b110111;     //123pi/512
   m_cos[123]  =  6'b001101;     //123pi/512
   m_sin[124]  =  6'b110111;     //124pi/512
   m_cos[124]  =  6'b001101;     //124pi/512
   m_sin[125]  =  6'b110111;     //125pi/512
   m_cos[125]  =  6'b001101;     //125pi/512
   m_sin[126]  =  6'b110111;     //126pi/512
   m_cos[126]  =  6'b001101;     //126pi/512
   m_sin[127]  =  6'b110111;     //127pi/512
   m_cos[127]  =  6'b001100;     //127pi/512
   m_sin[128]  =  6'b110111;     //128pi/512
   m_cos[128]  =  6'b001100;     //128pi/512
   m_sin[129]  =  6'b110111;     //129pi/512
   m_cos[129]  =  6'b001100;     //129pi/512
   m_sin[130]  =  6'b110110;     //130pi/512
   m_cos[130]  =  6'b001100;     //130pi/512
   m_sin[131]  =  6'b110110;     //131pi/512
   m_cos[131]  =  6'b001100;     //131pi/512
   m_sin[132]  =  6'b110110;     //132pi/512
   m_cos[132]  =  6'b001100;     //132pi/512
   m_sin[133]  =  6'b110110;     //133pi/512
   m_cos[133]  =  6'b001100;     //133pi/512
   m_sin[134]  =  6'b110110;     //134pi/512
   m_cos[134]  =  6'b001100;     //134pi/512
   m_sin[135]  =  6'b110110;     //135pi/512
   m_cos[135]  =  6'b001100;     //135pi/512
   m_sin[136]  =  6'b110110;     //136pi/512
   m_cos[136]  =  6'b001100;     //136pi/512
   m_sin[137]  =  6'b110110;     //137pi/512
   m_cos[137]  =  6'b001100;     //137pi/512
   m_sin[138]  =  6'b110110;     //138pi/512
   m_cos[138]  =  6'b001100;     //138pi/512
   m_sin[139]  =  6'b110110;     //139pi/512
   m_cos[139]  =  6'b001100;     //139pi/512
   m_sin[140]  =  6'b110110;     //140pi/512
   m_cos[140]  =  6'b001100;     //140pi/512
   m_sin[141]  =  6'b110110;     //141pi/512
   m_cos[141]  =  6'b001100;     //141pi/512
   m_sin[142]  =  6'b110110;     //142pi/512
   m_cos[142]  =  6'b001100;     //142pi/512
   m_sin[143]  =  6'b110110;     //143pi/512
   m_cos[143]  =  6'b001100;     //143pi/512
   m_sin[144]  =  6'b110110;     //144pi/512
   m_cos[144]  =  6'b001100;     //144pi/512
   m_sin[145]  =  6'b110110;     //145pi/512
   m_cos[145]  =  6'b001100;     //145pi/512
   m_sin[146]  =  6'b110101;     //146pi/512
   m_cos[146]  =  6'b001100;     //146pi/512
   m_sin[147]  =  6'b110101;     //147pi/512
   m_cos[147]  =  6'b001100;     //147pi/512
   m_sin[148]  =  6'b110101;     //148pi/512
   m_cos[148]  =  6'b001011;     //148pi/512
   m_sin[149]  =  6'b110101;     //149pi/512
   m_cos[149]  =  6'b001011;     //149pi/512
   m_sin[150]  =  6'b110101;     //150pi/512
   m_cos[150]  =  6'b001011;     //150pi/512
   m_sin[151]  =  6'b110101;     //151pi/512
   m_cos[151]  =  6'b001011;     //151pi/512
   m_sin[152]  =  6'b110101;     //152pi/512
   m_cos[152]  =  6'b001011;     //152pi/512
   m_sin[153]  =  6'b110101;     //153pi/512
   m_cos[153]  =  6'b001011;     //153pi/512
   m_sin[154]  =  6'b110101;     //154pi/512
   m_cos[154]  =  6'b001011;     //154pi/512
   m_sin[155]  =  6'b110101;     //155pi/512
   m_cos[155]  =  6'b001011;     //155pi/512
   m_sin[156]  =  6'b110101;     //156pi/512
   m_cos[156]  =  6'b001011;     //156pi/512
   m_sin[157]  =  6'b110101;     //157pi/512
   m_cos[157]  =  6'b001011;     //157pi/512
   m_sin[158]  =  6'b110101;     //158pi/512
   m_cos[158]  =  6'b001011;     //158pi/512
   m_sin[159]  =  6'b110101;     //159pi/512
   m_cos[159]  =  6'b001011;     //159pi/512
   m_sin[160]  =  6'b110101;     //160pi/512
   m_cos[160]  =  6'b001011;     //160pi/512
   m_sin[161]  =  6'b110101;     //161pi/512
   m_cos[161]  =  6'b001011;     //161pi/512
   m_sin[162]  =  6'b110101;     //162pi/512
   m_cos[162]  =  6'b001011;     //162pi/512
   m_sin[163]  =  6'b110101;     //163pi/512
   m_cos[163]  =  6'b001011;     //163pi/512
   m_sin[164]  =  6'b110100;     //164pi/512
   m_cos[164]  =  6'b001011;     //164pi/512
   m_sin[165]  =  6'b110100;     //165pi/512
   m_cos[165]  =  6'b001011;     //165pi/512
   m_sin[166]  =  6'b110100;     //166pi/512
   m_cos[166]  =  6'b001010;     //166pi/512
   m_sin[167]  =  6'b110100;     //167pi/512
   m_cos[167]  =  6'b001010;     //167pi/512
   m_sin[168]  =  6'b110100;     //168pi/512
   m_cos[168]  =  6'b001010;     //168pi/512
   m_sin[169]  =  6'b110100;     //169pi/512
   m_cos[169]  =  6'b001010;     //169pi/512
   m_sin[170]  =  6'b110100;     //170pi/512
   m_cos[170]  =  6'b001010;     //170pi/512
   m_sin[171]  =  6'b110100;     //171pi/512
   m_cos[171]  =  6'b001010;     //171pi/512
   m_sin[172]  =  6'b110100;     //172pi/512
   m_cos[172]  =  6'b001010;     //172pi/512
   m_sin[173]  =  6'b110100;     //173pi/512
   m_cos[173]  =  6'b001010;     //173pi/512
   m_sin[174]  =  6'b110100;     //174pi/512
   m_cos[174]  =  6'b001010;     //174pi/512
   m_sin[175]  =  6'b110100;     //175pi/512
   m_cos[175]  =  6'b001010;     //175pi/512
   m_sin[176]  =  6'b110100;     //176pi/512
   m_cos[176]  =  6'b001010;     //176pi/512
   m_sin[177]  =  6'b110100;     //177pi/512
   m_cos[177]  =  6'b001010;     //177pi/512
   m_sin[178]  =  6'b110100;     //178pi/512
   m_cos[178]  =  6'b001010;     //178pi/512
   m_sin[179]  =  6'b110100;     //179pi/512
   m_cos[179]  =  6'b001010;     //179pi/512
   m_sin[180]  =  6'b110100;     //180pi/512
   m_cos[180]  =  6'b001010;     //180pi/512
   m_sin[181]  =  6'b110100;     //181pi/512
   m_cos[181]  =  6'b001010;     //181pi/512
   m_sin[182]  =  6'b110100;     //182pi/512
   m_cos[182]  =  6'b001010;     //182pi/512
   m_sin[183]  =  6'b110011;     //183pi/512
   m_cos[183]  =  6'b001001;     //183pi/512
   m_sin[184]  =  6'b110011;     //184pi/512
   m_cos[184]  =  6'b001001;     //184pi/512
   m_sin[185]  =  6'b110011;     //185pi/512
   m_cos[185]  =  6'b001001;     //185pi/512
   m_sin[186]  =  6'b110011;     //186pi/512
   m_cos[186]  =  6'b001001;     //186pi/512
   m_sin[187]  =  6'b110011;     //187pi/512
   m_cos[187]  =  6'b001001;     //187pi/512
   m_sin[188]  =  6'b110011;     //188pi/512
   m_cos[188]  =  6'b001001;     //188pi/512
   m_sin[189]  =  6'b110011;     //189pi/512
   m_cos[189]  =  6'b001001;     //189pi/512
   m_sin[190]  =  6'b110011;     //190pi/512
   m_cos[190]  =  6'b001001;     //190pi/512
   m_sin[191]  =  6'b110011;     //191pi/512
   m_cos[191]  =  6'b001001;     //191pi/512
   m_sin[192]  =  6'b110011;     //192pi/512
   m_cos[192]  =  6'b001001;     //192pi/512
   m_sin[193]  =  6'b110011;     //193pi/512
   m_cos[193]  =  6'b001001;     //193pi/512
   m_sin[194]  =  6'b110011;     //194pi/512
   m_cos[194]  =  6'b001001;     //194pi/512
   m_sin[195]  =  6'b110011;     //195pi/512
   m_cos[195]  =  6'b001001;     //195pi/512
   m_sin[196]  =  6'b110011;     //196pi/512
   m_cos[196]  =  6'b001001;     //196pi/512
   m_sin[197]  =  6'b110011;     //197pi/512
   m_cos[197]  =  6'b001001;     //197pi/512
   m_sin[198]  =  6'b110011;     //198pi/512
   m_cos[198]  =  6'b001001;     //198pi/512
   m_sin[199]  =  6'b110011;     //199pi/512
   m_cos[199]  =  6'b001000;     //199pi/512
   m_sin[200]  =  6'b110011;     //200pi/512
   m_cos[200]  =  6'b001000;     //200pi/512
   m_sin[201]  =  6'b110011;     //201pi/512
   m_cos[201]  =  6'b001000;     //201pi/512
   m_sin[202]  =  6'b110011;     //202pi/512
   m_cos[202]  =  6'b001000;     //202pi/512
   m_sin[203]  =  6'b110011;     //203pi/512
   m_cos[203]  =  6'b001000;     //203pi/512
   m_sin[204]  =  6'b110011;     //204pi/512
   m_cos[204]  =  6'b001000;     //204pi/512
   m_sin[205]  =  6'b110010;     //205pi/512
   m_cos[205]  =  6'b001000;     //205pi/512
   m_sin[206]  =  6'b110010;     //206pi/512
   m_cos[206]  =  6'b001000;     //206pi/512
   m_sin[207]  =  6'b110010;     //207pi/512
   m_cos[207]  =  6'b001000;     //207pi/512
   m_sin[208]  =  6'b110010;     //208pi/512
   m_cos[208]  =  6'b001000;     //208pi/512
   m_sin[209]  =  6'b110010;     //209pi/512
   m_cos[209]  =  6'b001000;     //209pi/512
   m_sin[210]  =  6'b110010;     //210pi/512
   m_cos[210]  =  6'b001000;     //210pi/512
   m_sin[211]  =  6'b110010;     //211pi/512
   m_cos[211]  =  6'b001000;     //211pi/512
   m_sin[212]  =  6'b110010;     //212pi/512
   m_cos[212]  =  6'b001000;     //212pi/512
   m_sin[213]  =  6'b110010;     //213pi/512
   m_cos[213]  =  6'b001000;     //213pi/512
   m_sin[214]  =  6'b110010;     //214pi/512
   m_cos[214]  =  6'b000111;     //214pi/512
   m_sin[215]  =  6'b110010;     //215pi/512
   m_cos[215]  =  6'b000111;     //215pi/512
   m_sin[216]  =  6'b110010;     //216pi/512
   m_cos[216]  =  6'b000111;     //216pi/512
   m_sin[217]  =  6'b110010;     //217pi/512
   m_cos[217]  =  6'b000111;     //217pi/512
   m_sin[218]  =  6'b110010;     //218pi/512
   m_cos[218]  =  6'b000111;     //218pi/512
   m_sin[219]  =  6'b110010;     //219pi/512
   m_cos[219]  =  6'b000111;     //219pi/512
   m_sin[220]  =  6'b110010;     //220pi/512
   m_cos[220]  =  6'b000111;     //220pi/512
   m_sin[221]  =  6'b110010;     //221pi/512
   m_cos[221]  =  6'b000111;     //221pi/512
   m_sin[222]  =  6'b110010;     //222pi/512
   m_cos[222]  =  6'b000111;     //222pi/512
   m_sin[223]  =  6'b110010;     //223pi/512
   m_cos[223]  =  6'b000111;     //223pi/512
   m_sin[224]  =  6'b110010;     //224pi/512
   m_cos[224]  =  6'b000111;     //224pi/512
   m_sin[225]  =  6'b110010;     //225pi/512
   m_cos[225]  =  6'b000111;     //225pi/512
   m_sin[226]  =  6'b110010;     //226pi/512
   m_cos[226]  =  6'b000111;     //226pi/512
   m_sin[227]  =  6'b110010;     //227pi/512
   m_cos[227]  =  6'b000111;     //227pi/512
   m_sin[228]  =  6'b110010;     //228pi/512
   m_cos[228]  =  6'b000110;     //228pi/512
   m_sin[229]  =  6'b110010;     //229pi/512
   m_cos[229]  =  6'b000110;     //229pi/512
   m_sin[230]  =  6'b110010;     //230pi/512
   m_cos[230]  =  6'b000110;     //230pi/512
   m_sin[231]  =  6'b110010;     //231pi/512
   m_cos[231]  =  6'b000110;     //231pi/512
   m_sin[232]  =  6'b110001;     //232pi/512
   m_cos[232]  =  6'b000110;     //232pi/512
   m_sin[233]  =  6'b110001;     //233pi/512
   m_cos[233]  =  6'b000110;     //233pi/512
   m_sin[234]  =  6'b110001;     //234pi/512
   m_cos[234]  =  6'b000110;     //234pi/512
   m_sin[235]  =  6'b110001;     //235pi/512
   m_cos[235]  =  6'b000110;     //235pi/512
   m_sin[236]  =  6'b110001;     //236pi/512
   m_cos[236]  =  6'b000110;     //236pi/512
   m_sin[237]  =  6'b110001;     //237pi/512
   m_cos[237]  =  6'b000110;     //237pi/512
   m_sin[238]  =  6'b110001;     //238pi/512
   m_cos[238]  =  6'b000110;     //238pi/512
   m_sin[239]  =  6'b110001;     //239pi/512
   m_cos[239]  =  6'b000110;     //239pi/512
   m_sin[240]  =  6'b110001;     //240pi/512
   m_cos[240]  =  6'b000110;     //240pi/512
   m_sin[241]  =  6'b110001;     //241pi/512
   m_cos[241]  =  6'b000110;     //241pi/512
   m_sin[242]  =  6'b110001;     //242pi/512
   m_cos[242]  =  6'b000101;     //242pi/512
   m_sin[243]  =  6'b110001;     //243pi/512
   m_cos[243]  =  6'b000101;     //243pi/512
   m_sin[244]  =  6'b110001;     //244pi/512
   m_cos[244]  =  6'b000101;     //244pi/512
   m_sin[245]  =  6'b110001;     //245pi/512
   m_cos[245]  =  6'b000101;     //245pi/512
   m_sin[246]  =  6'b110001;     //246pi/512
   m_cos[246]  =  6'b000101;     //246pi/512
   m_sin[247]  =  6'b110001;     //247pi/512
   m_cos[247]  =  6'b000101;     //247pi/512
   m_sin[248]  =  6'b110001;     //248pi/512
   m_cos[248]  =  6'b000101;     //248pi/512
   m_sin[249]  =  6'b110001;     //249pi/512
   m_cos[249]  =  6'b000101;     //249pi/512
   m_sin[250]  =  6'b110001;     //250pi/512
   m_cos[250]  =  6'b000101;     //250pi/512
   m_sin[251]  =  6'b110001;     //251pi/512
   m_cos[251]  =  6'b000101;     //251pi/512
   m_sin[252]  =  6'b110001;     //252pi/512
   m_cos[252]  =  6'b000101;     //252pi/512
   m_sin[253]  =  6'b110001;     //253pi/512
   m_cos[253]  =  6'b000101;     //253pi/512
   m_sin[254]  =  6'b110001;     //254pi/512
   m_cos[254]  =  6'b000101;     //254pi/512
   m_sin[255]  =  6'b110001;     //255pi/512
   m_cos[255]  =  6'b000101;     //255pi/512
   m_sin[256]  =  6'b110001;     //256pi/512
   m_cos[256]  =  6'b000100;     //256pi/512
   m_sin[257]  =  6'b110001;     //257pi/512
   m_cos[257]  =  6'b000100;     //257pi/512
   m_sin[258]  =  6'b110001;     //258pi/512
   m_cos[258]  =  6'b000100;     //258pi/512
   m_sin[259]  =  6'b110001;     //259pi/512
   m_cos[259]  =  6'b000100;     //259pi/512
   m_sin[260]  =  6'b110001;     //260pi/512
   m_cos[260]  =  6'b000100;     //260pi/512
   m_sin[261]  =  6'b110001;     //261pi/512
   m_cos[261]  =  6'b000100;     //261pi/512
   m_sin[262]  =  6'b110001;     //262pi/512
   m_cos[262]  =  6'b000100;     //262pi/512
   m_sin[263]  =  6'b110001;     //263pi/512
   m_cos[263]  =  6'b000100;     //263pi/512
   m_sin[264]  =  6'b110001;     //264pi/512
   m_cos[264]  =  6'b000100;     //264pi/512
   m_sin[265]  =  6'b110001;     //265pi/512
   m_cos[265]  =  6'b000100;     //265pi/512
   m_sin[266]  =  6'b110001;     //266pi/512
   m_cos[266]  =  6'b000100;     //266pi/512
   m_sin[267]  =  6'b110001;     //267pi/512
   m_cos[267]  =  6'b000100;     //267pi/512
   m_sin[268]  =  6'b110001;     //268pi/512
   m_cos[268]  =  6'b000100;     //268pi/512
   m_sin[269]  =  6'b110000;     //269pi/512
   m_cos[269]  =  6'b000011;     //269pi/512
   m_sin[270]  =  6'b110000;     //270pi/512
   m_cos[270]  =  6'b000011;     //270pi/512
   m_sin[271]  =  6'b110000;     //271pi/512
   m_cos[271]  =  6'b000011;     //271pi/512
   m_sin[272]  =  6'b110000;     //272pi/512
   m_cos[272]  =  6'b000011;     //272pi/512
   m_sin[273]  =  6'b110000;     //273pi/512
   m_cos[273]  =  6'b000011;     //273pi/512
   m_sin[274]  =  6'b110000;     //274pi/512
   m_cos[274]  =  6'b000011;     //274pi/512
   m_sin[275]  =  6'b110000;     //275pi/512
   m_cos[275]  =  6'b000011;     //275pi/512
   m_sin[276]  =  6'b110000;     //276pi/512
   m_cos[276]  =  6'b000011;     //276pi/512
   m_sin[277]  =  6'b110000;     //277pi/512
   m_cos[277]  =  6'b000011;     //277pi/512
   m_sin[278]  =  6'b110000;     //278pi/512
   m_cos[278]  =  6'b000011;     //278pi/512
   m_sin[279]  =  6'b110000;     //279pi/512
   m_cos[279]  =  6'b000011;     //279pi/512
   m_sin[280]  =  6'b110000;     //280pi/512
   m_cos[280]  =  6'b000011;     //280pi/512
   m_sin[281]  =  6'b110000;     //281pi/512
   m_cos[281]  =  6'b000011;     //281pi/512
   m_sin[282]  =  6'b110000;     //282pi/512
   m_cos[282]  =  6'b000010;     //282pi/512
   m_sin[283]  =  6'b110000;     //283pi/512
   m_cos[283]  =  6'b000010;     //283pi/512
   m_sin[284]  =  6'b110000;     //284pi/512
   m_cos[284]  =  6'b000010;     //284pi/512
   m_sin[285]  =  6'b110000;     //285pi/512
   m_cos[285]  =  6'b000010;     //285pi/512
   m_sin[286]  =  6'b110000;     //286pi/512
   m_cos[286]  =  6'b000010;     //286pi/512
   m_sin[287]  =  6'b110000;     //287pi/512
   m_cos[287]  =  6'b000010;     //287pi/512
   m_sin[288]  =  6'b110000;     //288pi/512
   m_cos[288]  =  6'b000010;     //288pi/512
   m_sin[289]  =  6'b110000;     //289pi/512
   m_cos[289]  =  6'b000010;     //289pi/512
   m_sin[290]  =  6'b110000;     //290pi/512
   m_cos[290]  =  6'b000010;     //290pi/512
   m_sin[291]  =  6'b110000;     //291pi/512
   m_cos[291]  =  6'b000010;     //291pi/512
   m_sin[292]  =  6'b110000;     //292pi/512
   m_cos[292]  =  6'b000010;     //292pi/512
   m_sin[293]  =  6'b110000;     //293pi/512
   m_cos[293]  =  6'b000010;     //293pi/512
   m_sin[294]  =  6'b110000;     //294pi/512
   m_cos[294]  =  6'b000010;     //294pi/512
   m_sin[295]  =  6'b110000;     //295pi/512
   m_cos[295]  =  6'b000001;     //295pi/512
   m_sin[296]  =  6'b110000;     //296pi/512
   m_cos[296]  =  6'b000001;     //296pi/512
   m_sin[297]  =  6'b110000;     //297pi/512
   m_cos[297]  =  6'b000001;     //297pi/512
   m_sin[298]  =  6'b110000;     //298pi/512
   m_cos[298]  =  6'b000001;     //298pi/512
   m_sin[299]  =  6'b110000;     //299pi/512
   m_cos[299]  =  6'b000001;     //299pi/512
   m_sin[300]  =  6'b110000;     //300pi/512
   m_cos[300]  =  6'b000001;     //300pi/512
   m_sin[301]  =  6'b110000;     //301pi/512
   m_cos[301]  =  6'b000001;     //301pi/512
   m_sin[302]  =  6'b110000;     //302pi/512
   m_cos[302]  =  6'b000001;     //302pi/512
   m_sin[303]  =  6'b110000;     //303pi/512
   m_cos[303]  =  6'b000001;     //303pi/512
   m_sin[304]  =  6'b110000;     //304pi/512
   m_cos[304]  =  6'b000001;     //304pi/512
   m_sin[305]  =  6'b110000;     //305pi/512
   m_cos[305]  =  6'b000001;     //305pi/512
   m_sin[306]  =  6'b110000;     //306pi/512
   m_cos[306]  =  6'b000001;     //306pi/512
   m_sin[307]  =  6'b110000;     //307pi/512
   m_cos[307]  =  6'b000001;     //307pi/512
   m_sin[308]  =  6'b110000;     //308pi/512
   m_cos[308]  =  6'b000000;     //308pi/512
   m_sin[309]  =  6'b110000;     //309pi/512
   m_cos[309]  =  6'b000000;     //309pi/512
   m_sin[310]  =  6'b110000;     //310pi/512
   m_cos[310]  =  6'b000000;     //310pi/512
   m_sin[311]  =  6'b110000;     //311pi/512
   m_cos[311]  =  6'b000000;     //311pi/512
   m_sin[312]  =  6'b110000;     //312pi/512
   m_cos[312]  =  6'b000000;     //312pi/512
   m_sin[313]  =  6'b110000;     //313pi/512
   m_cos[313]  =  6'b000000;     //313pi/512
   m_sin[314]  =  6'b110000;     //314pi/512
   m_cos[314]  =  6'b000000;     //314pi/512
   m_sin[315]  =  6'b110000;     //315pi/512
   m_cos[315]  =  6'b000000;     //315pi/512
   m_sin[316]  =  6'b110000;     //316pi/512
   m_cos[316]  =  6'b000000;     //316pi/512
   m_sin[317]  =  6'b110000;     //317pi/512
   m_cos[317]  =  6'b000000;     //317pi/512
   m_sin[318]  =  6'b110000;     //318pi/512
   m_cos[318]  =  6'b000000;     //318pi/512
   m_sin[319]  =  6'b110000;     //319pi/512
   m_cos[319]  =  6'b000000;     //319pi/512
   m_sin[320]  =  6'b110000;     //320pi/512
   m_cos[320]  =  6'b000000;     //320pi/512
   m_sin[321]  =  6'b110000;     //321pi/512
   m_cos[321]  =  6'b000000;     //321pi/512
   m_sin[322]  =  6'b110000;     //322pi/512
   m_cos[322]  =  6'b000000;     //322pi/512
   m_sin[323]  =  6'b110000;     //323pi/512
   m_cos[323]  =  6'b000000;     //323pi/512
   m_sin[324]  =  6'b110000;     //324pi/512
   m_cos[324]  =  6'b000000;     //324pi/512
   m_sin[325]  =  6'b110000;     //325pi/512
   m_cos[325]  =  6'b000000;     //325pi/512
   m_sin[326]  =  6'b110000;     //326pi/512
   m_cos[326]  =  6'b000000;     //326pi/512
   m_sin[327]  =  6'b110000;     //327pi/512
   m_cos[327]  =  6'b111111;     //327pi/512
   m_sin[328]  =  6'b110000;     //328pi/512
   m_cos[328]  =  6'b111111;     //328pi/512
   m_sin[329]  =  6'b110000;     //329pi/512
   m_cos[329]  =  6'b111111;     //329pi/512
   m_sin[330]  =  6'b110000;     //330pi/512
   m_cos[330]  =  6'b111111;     //330pi/512
   m_sin[331]  =  6'b110000;     //331pi/512
   m_cos[331]  =  6'b111111;     //331pi/512
   m_sin[332]  =  6'b110000;     //332pi/512
   m_cos[332]  =  6'b111111;     //332pi/512
   m_sin[333]  =  6'b110000;     //333pi/512
   m_cos[333]  =  6'b111111;     //333pi/512
   m_sin[334]  =  6'b110000;     //334pi/512
   m_cos[334]  =  6'b111111;     //334pi/512
   m_sin[335]  =  6'b110000;     //335pi/512
   m_cos[335]  =  6'b111111;     //335pi/512
   m_sin[336]  =  6'b110000;     //336pi/512
   m_cos[336]  =  6'b111111;     //336pi/512
   m_sin[337]  =  6'b110000;     //337pi/512
   m_cos[337]  =  6'b111111;     //337pi/512
   m_sin[338]  =  6'b110000;     //338pi/512
   m_cos[338]  =  6'b111111;     //338pi/512
   m_sin[339]  =  6'b110000;     //339pi/512
   m_cos[339]  =  6'b111111;     //339pi/512
   m_sin[340]  =  6'b110000;     //340pi/512
   m_cos[340]  =  6'b111110;     //340pi/512
   m_sin[341]  =  6'b110000;     //341pi/512
   m_cos[341]  =  6'b111110;     //341pi/512
   m_sin[342]  =  6'b110000;     //342pi/512
   m_cos[342]  =  6'b111110;     //342pi/512
   m_sin[343]  =  6'b110000;     //343pi/512
   m_cos[343]  =  6'b111110;     //343pi/512
   m_sin[344]  =  6'b110000;     //344pi/512
   m_cos[344]  =  6'b111110;     //344pi/512
   m_sin[345]  =  6'b110000;     //345pi/512
   m_cos[345]  =  6'b111110;     //345pi/512
   m_sin[346]  =  6'b110000;     //346pi/512
   m_cos[346]  =  6'b111110;     //346pi/512
   m_sin[347]  =  6'b110000;     //347pi/512
   m_cos[347]  =  6'b111110;     //347pi/512
   m_sin[348]  =  6'b110000;     //348pi/512
   m_cos[348]  =  6'b111110;     //348pi/512
   m_sin[349]  =  6'b110000;     //349pi/512
   m_cos[349]  =  6'b111110;     //349pi/512
   m_sin[350]  =  6'b110000;     //350pi/512
   m_cos[350]  =  6'b111110;     //350pi/512
   m_sin[351]  =  6'b110000;     //351pi/512
   m_cos[351]  =  6'b111110;     //351pi/512
   m_sin[352]  =  6'b110000;     //352pi/512
   m_cos[352]  =  6'b111101;     //352pi/512
   m_sin[353]  =  6'b110000;     //353pi/512
   m_cos[353]  =  6'b111101;     //353pi/512
   m_sin[354]  =  6'b110000;     //354pi/512
   m_cos[354]  =  6'b111101;     //354pi/512
   m_sin[355]  =  6'b110000;     //355pi/512
   m_cos[355]  =  6'b111101;     //355pi/512
   m_sin[356]  =  6'b110000;     //356pi/512
   m_cos[356]  =  6'b111101;     //356pi/512
   m_sin[357]  =  6'b110000;     //357pi/512
   m_cos[357]  =  6'b111101;     //357pi/512
   m_sin[358]  =  6'b110000;     //358pi/512
   m_cos[358]  =  6'b111101;     //358pi/512
   m_sin[359]  =  6'b110000;     //359pi/512
   m_cos[359]  =  6'b111101;     //359pi/512
   m_sin[360]  =  6'b110000;     //360pi/512
   m_cos[360]  =  6'b111101;     //360pi/512
   m_sin[361]  =  6'b110000;     //361pi/512
   m_cos[361]  =  6'b111101;     //361pi/512
   m_sin[362]  =  6'b110000;     //362pi/512
   m_cos[362]  =  6'b111101;     //362pi/512
   m_sin[363]  =  6'b110000;     //363pi/512
   m_cos[363]  =  6'b111101;     //363pi/512
   m_sin[364]  =  6'b110000;     //364pi/512
   m_cos[364]  =  6'b111101;     //364pi/512
   m_sin[365]  =  6'b110000;     //365pi/512
   m_cos[365]  =  6'b111100;     //365pi/512
   m_sin[366]  =  6'b110000;     //366pi/512
   m_cos[366]  =  6'b111100;     //366pi/512
   m_sin[367]  =  6'b110000;     //367pi/512
   m_cos[367]  =  6'b111100;     //367pi/512
   m_sin[368]  =  6'b110000;     //368pi/512
   m_cos[368]  =  6'b111100;     //368pi/512
   m_sin[369]  =  6'b110000;     //369pi/512
   m_cos[369]  =  6'b111100;     //369pi/512
   m_sin[370]  =  6'b110000;     //370pi/512
   m_cos[370]  =  6'b111100;     //370pi/512
   m_sin[371]  =  6'b110000;     //371pi/512
   m_cos[371]  =  6'b111100;     //371pi/512
   m_sin[372]  =  6'b110001;     //372pi/512
   m_cos[372]  =  6'b111100;     //372pi/512
   m_sin[373]  =  6'b110001;     //373pi/512
   m_cos[373]  =  6'b111100;     //373pi/512
   m_sin[374]  =  6'b110001;     //374pi/512
   m_cos[374]  =  6'b111100;     //374pi/512
   m_sin[375]  =  6'b110001;     //375pi/512
   m_cos[375]  =  6'b111100;     //375pi/512
   m_sin[376]  =  6'b110001;     //376pi/512
   m_cos[376]  =  6'b111100;     //376pi/512
   m_sin[377]  =  6'b110001;     //377pi/512
   m_cos[377]  =  6'b111100;     //377pi/512
   m_sin[378]  =  6'b110001;     //378pi/512
   m_cos[378]  =  6'b111100;     //378pi/512
   m_sin[379]  =  6'b110001;     //379pi/512
   m_cos[379]  =  6'b111011;     //379pi/512
   m_sin[380]  =  6'b110001;     //380pi/512
   m_cos[380]  =  6'b111011;     //380pi/512
   m_sin[381]  =  6'b110001;     //381pi/512
   m_cos[381]  =  6'b111011;     //381pi/512
   m_sin[382]  =  6'b110001;     //382pi/512
   m_cos[382]  =  6'b111011;     //382pi/512
   m_sin[383]  =  6'b110001;     //383pi/512
   m_cos[383]  =  6'b111011;     //383pi/512
   m_sin[384]  =  6'b110001;     //384pi/512
   m_cos[384]  =  6'b111011;     //384pi/512
   m_sin[385]  =  6'b110001;     //385pi/512
   m_cos[385]  =  6'b111011;     //385pi/512
   m_sin[386]  =  6'b110001;     //386pi/512
   m_cos[386]  =  6'b111011;     //386pi/512
   m_sin[387]  =  6'b110001;     //387pi/512
   m_cos[387]  =  6'b111011;     //387pi/512
   m_sin[388]  =  6'b110001;     //388pi/512
   m_cos[388]  =  6'b111011;     //388pi/512
   m_sin[389]  =  6'b110001;     //389pi/512
   m_cos[389]  =  6'b111011;     //389pi/512
   m_sin[390]  =  6'b110001;     //390pi/512
   m_cos[390]  =  6'b111011;     //390pi/512
   m_sin[391]  =  6'b110001;     //391pi/512
   m_cos[391]  =  6'b111011;     //391pi/512
   m_sin[392]  =  6'b110001;     //392pi/512
   m_cos[392]  =  6'b111010;     //392pi/512
   m_sin[393]  =  6'b110001;     //393pi/512
   m_cos[393]  =  6'b111010;     //393pi/512
   m_sin[394]  =  6'b110001;     //394pi/512
   m_cos[394]  =  6'b111010;     //394pi/512
   m_sin[395]  =  6'b110001;     //395pi/512
   m_cos[395]  =  6'b111010;     //395pi/512
   m_sin[396]  =  6'b110001;     //396pi/512
   m_cos[396]  =  6'b111010;     //396pi/512
   m_sin[397]  =  6'b110001;     //397pi/512
   m_cos[397]  =  6'b111010;     //397pi/512
   m_sin[398]  =  6'b110001;     //398pi/512
   m_cos[398]  =  6'b111010;     //398pi/512
   m_sin[399]  =  6'b110001;     //399pi/512
   m_cos[399]  =  6'b111010;     //399pi/512
   m_sin[400]  =  6'b110001;     //400pi/512
   m_cos[400]  =  6'b111010;     //400pi/512
   m_sin[401]  =  6'b110001;     //401pi/512
   m_cos[401]  =  6'b111010;     //401pi/512
   m_sin[402]  =  6'b110001;     //402pi/512
   m_cos[402]  =  6'b111010;     //402pi/512
   m_sin[403]  =  6'b110001;     //403pi/512
   m_cos[403]  =  6'b111010;     //403pi/512
   m_sin[404]  =  6'b110001;     //404pi/512
   m_cos[404]  =  6'b111010;     //404pi/512
   m_sin[405]  =  6'b110001;     //405pi/512
   m_cos[405]  =  6'b111010;     //405pi/512
   m_sin[406]  =  6'b110001;     //406pi/512
   m_cos[406]  =  6'b111001;     //406pi/512
   m_sin[407]  =  6'b110001;     //407pi/512
   m_cos[407]  =  6'b111001;     //407pi/512
   m_sin[408]  =  6'b110001;     //408pi/512
   m_cos[408]  =  6'b111001;     //408pi/512
   m_sin[409]  =  6'b110010;     //409pi/512
   m_cos[409]  =  6'b111001;     //409pi/512
   m_sin[410]  =  6'b110010;     //410pi/512
   m_cos[410]  =  6'b111001;     //410pi/512
   m_sin[411]  =  6'b110010;     //411pi/512
   m_cos[411]  =  6'b111001;     //411pi/512
   m_sin[412]  =  6'b110010;     //412pi/512
   m_cos[412]  =  6'b111001;     //412pi/512
   m_sin[413]  =  6'b110010;     //413pi/512
   m_cos[413]  =  6'b111001;     //413pi/512
   m_sin[414]  =  6'b110010;     //414pi/512
   m_cos[414]  =  6'b111001;     //414pi/512
   m_sin[415]  =  6'b110010;     //415pi/512
   m_cos[415]  =  6'b111001;     //415pi/512
   m_sin[416]  =  6'b110010;     //416pi/512
   m_cos[416]  =  6'b111001;     //416pi/512
   m_sin[417]  =  6'b110010;     //417pi/512
   m_cos[417]  =  6'b111001;     //417pi/512
   m_sin[418]  =  6'b110010;     //418pi/512
   m_cos[418]  =  6'b111001;     //418pi/512
   m_sin[419]  =  6'b110010;     //419pi/512
   m_cos[419]  =  6'b111001;     //419pi/512
   m_sin[420]  =  6'b110010;     //420pi/512
   m_cos[420]  =  6'b111000;     //420pi/512
   m_sin[421]  =  6'b110010;     //421pi/512
   m_cos[421]  =  6'b111000;     //421pi/512
   m_sin[422]  =  6'b110010;     //422pi/512
   m_cos[422]  =  6'b111000;     //422pi/512
   m_sin[423]  =  6'b110010;     //423pi/512
   m_cos[423]  =  6'b111000;     //423pi/512
   m_sin[424]  =  6'b110010;     //424pi/512
   m_cos[424]  =  6'b111000;     //424pi/512
   m_sin[425]  =  6'b110010;     //425pi/512
   m_cos[425]  =  6'b111000;     //425pi/512
   m_sin[426]  =  6'b110010;     //426pi/512
   m_cos[426]  =  6'b111000;     //426pi/512
   m_sin[427]  =  6'b110010;     //427pi/512
   m_cos[427]  =  6'b111000;     //427pi/512
   m_sin[428]  =  6'b110010;     //428pi/512
   m_cos[428]  =  6'b111000;     //428pi/512
   m_sin[429]  =  6'b110010;     //429pi/512
   m_cos[429]  =  6'b111000;     //429pi/512
   m_sin[430]  =  6'b110010;     //430pi/512
   m_cos[430]  =  6'b111000;     //430pi/512
   m_sin[431]  =  6'b110010;     //431pi/512
   m_cos[431]  =  6'b111000;     //431pi/512
   m_sin[432]  =  6'b110010;     //432pi/512
   m_cos[432]  =  6'b111000;     //432pi/512
   m_sin[433]  =  6'b110010;     //433pi/512
   m_cos[433]  =  6'b111000;     //433pi/512
   m_sin[434]  =  6'b110010;     //434pi/512
   m_cos[434]  =  6'b111000;     //434pi/512
   m_sin[435]  =  6'b110010;     //435pi/512
   m_cos[435]  =  6'b110111;     //435pi/512
   m_sin[436]  =  6'b110011;     //436pi/512
   m_cos[436]  =  6'b110111;     //436pi/512
   m_sin[437]  =  6'b110011;     //437pi/512
   m_cos[437]  =  6'b110111;     //437pi/512
   m_sin[438]  =  6'b110011;     //438pi/512
   m_cos[438]  =  6'b110111;     //438pi/512
   m_sin[439]  =  6'b110011;     //439pi/512
   m_cos[439]  =  6'b110111;     //439pi/512
   m_sin[440]  =  6'b110011;     //440pi/512
   m_cos[440]  =  6'b110111;     //440pi/512
   m_sin[441]  =  6'b110011;     //441pi/512
   m_cos[441]  =  6'b110111;     //441pi/512
   m_sin[442]  =  6'b110011;     //442pi/512
   m_cos[442]  =  6'b110111;     //442pi/512
   m_sin[443]  =  6'b110011;     //443pi/512
   m_cos[443]  =  6'b110111;     //443pi/512
   m_sin[444]  =  6'b110011;     //444pi/512
   m_cos[444]  =  6'b110111;     //444pi/512
   m_sin[445]  =  6'b110011;     //445pi/512
   m_cos[445]  =  6'b110111;     //445pi/512
   m_sin[446]  =  6'b110011;     //446pi/512
   m_cos[446]  =  6'b110111;     //446pi/512
   m_sin[447]  =  6'b110011;     //447pi/512
   m_cos[447]  =  6'b110111;     //447pi/512
   m_sin[448]  =  6'b110011;     //448pi/512
   m_cos[448]  =  6'b110111;     //448pi/512
   m_sin[449]  =  6'b110011;     //449pi/512
   m_cos[449]  =  6'b110111;     //449pi/512
   m_sin[450]  =  6'b110011;     //450pi/512
   m_cos[450]  =  6'b110110;     //450pi/512
   m_sin[451]  =  6'b110011;     //451pi/512
   m_cos[451]  =  6'b110110;     //451pi/512
   m_sin[452]  =  6'b110011;     //452pi/512
   m_cos[452]  =  6'b110110;     //452pi/512
   m_sin[453]  =  6'b110011;     //453pi/512
   m_cos[453]  =  6'b110110;     //453pi/512
   m_sin[454]  =  6'b110011;     //454pi/512
   m_cos[454]  =  6'b110110;     //454pi/512
   m_sin[455]  =  6'b110011;     //455pi/512
   m_cos[455]  =  6'b110110;     //455pi/512
   m_sin[456]  =  6'b110011;     //456pi/512
   m_cos[456]  =  6'b110110;     //456pi/512
   m_sin[457]  =  6'b110011;     //457pi/512
   m_cos[457]  =  6'b110110;     //457pi/512
   m_sin[458]  =  6'b110100;     //458pi/512
   m_cos[458]  =  6'b110110;     //458pi/512
   m_sin[459]  =  6'b110100;     //459pi/512
   m_cos[459]  =  6'b110110;     //459pi/512
   m_sin[460]  =  6'b110100;     //460pi/512
   m_cos[460]  =  6'b110110;     //460pi/512
   m_sin[461]  =  6'b110100;     //461pi/512
   m_cos[461]  =  6'b110110;     //461pi/512
   m_sin[462]  =  6'b110100;     //462pi/512
   m_cos[462]  =  6'b110110;     //462pi/512
   m_sin[463]  =  6'b110100;     //463pi/512
   m_cos[463]  =  6'b110110;     //463pi/512
   m_sin[464]  =  6'b110100;     //464pi/512
   m_cos[464]  =  6'b110110;     //464pi/512
   m_sin[465]  =  6'b110100;     //465pi/512
   m_cos[465]  =  6'b110110;     //465pi/512
   m_sin[466]  =  6'b110100;     //466pi/512
   m_cos[466]  =  6'b110101;     //466pi/512
   m_sin[467]  =  6'b110100;     //467pi/512
   m_cos[467]  =  6'b110101;     //467pi/512
   m_sin[468]  =  6'b110100;     //468pi/512
   m_cos[468]  =  6'b110101;     //468pi/512
   m_sin[469]  =  6'b110100;     //469pi/512
   m_cos[469]  =  6'b110101;     //469pi/512
   m_sin[470]  =  6'b110100;     //470pi/512
   m_cos[470]  =  6'b110101;     //470pi/512
   m_sin[471]  =  6'b110100;     //471pi/512
   m_cos[471]  =  6'b110101;     //471pi/512
   m_sin[472]  =  6'b110100;     //472pi/512
   m_cos[472]  =  6'b110101;     //472pi/512
   m_sin[473]  =  6'b110100;     //473pi/512
   m_cos[473]  =  6'b110101;     //473pi/512
   m_sin[474]  =  6'b110100;     //474pi/512
   m_cos[474]  =  6'b110101;     //474pi/512
   m_sin[475]  =  6'b110100;     //475pi/512
   m_cos[475]  =  6'b110101;     //475pi/512
   m_sin[476]  =  6'b110100;     //476pi/512
   m_cos[476]  =  6'b110101;     //476pi/512
   m_sin[477]  =  6'b110101;     //477pi/512
   m_cos[477]  =  6'b110101;     //477pi/512
   m_sin[478]  =  6'b110101;     //478pi/512
   m_cos[478]  =  6'b110101;     //478pi/512
   m_sin[479]  =  6'b110101;     //479pi/512
   m_cos[479]  =  6'b110101;     //479pi/512
   m_sin[480]  =  6'b110101;     //480pi/512
   m_cos[480]  =  6'b110101;     //480pi/512
   m_sin[481]  =  6'b110101;     //481pi/512
   m_cos[481]  =  6'b110101;     //481pi/512
   m_sin[482]  =  6'b110101;     //482pi/512
   m_cos[482]  =  6'b110101;     //482pi/512
   m_sin[483]  =  6'b110101;     //483pi/512
   m_cos[483]  =  6'b110101;     //483pi/512
   m_sin[484]  =  6'b110101;     //484pi/512
   m_cos[484]  =  6'b110100;     //484pi/512
   m_sin[485]  =  6'b110101;     //485pi/512
   m_cos[485]  =  6'b110100;     //485pi/512
   m_sin[486]  =  6'b110101;     //486pi/512
   m_cos[486]  =  6'b110100;     //486pi/512
   m_sin[487]  =  6'b110101;     //487pi/512
   m_cos[487]  =  6'b110100;     //487pi/512
   m_sin[488]  =  6'b110101;     //488pi/512
   m_cos[488]  =  6'b110100;     //488pi/512
   m_sin[489]  =  6'b110101;     //489pi/512
   m_cos[489]  =  6'b110100;     //489pi/512
   m_sin[490]  =  6'b110101;     //490pi/512
   m_cos[490]  =  6'b110100;     //490pi/512
   m_sin[491]  =  6'b110101;     //491pi/512
   m_cos[491]  =  6'b110100;     //491pi/512
   m_sin[492]  =  6'b110101;     //492pi/512
   m_cos[492]  =  6'b110100;     //492pi/512
   m_sin[493]  =  6'b110101;     //493pi/512
   m_cos[493]  =  6'b110100;     //493pi/512
   m_sin[494]  =  6'b110101;     //494pi/512
   m_cos[494]  =  6'b110100;     //494pi/512
   m_sin[495]  =  6'b110110;     //495pi/512
   m_cos[495]  =  6'b110100;     //495pi/512
   m_sin[496]  =  6'b110110;     //496pi/512
   m_cos[496]  =  6'b110100;     //496pi/512
   m_sin[497]  =  6'b110110;     //497pi/512
   m_cos[497]  =  6'b110100;     //497pi/512
   m_sin[498]  =  6'b110110;     //498pi/512
   m_cos[498]  =  6'b110100;     //498pi/512
   m_sin[499]  =  6'b110110;     //499pi/512
   m_cos[499]  =  6'b110100;     //499pi/512
   m_sin[500]  =  6'b110110;     //500pi/512
   m_cos[500]  =  6'b110100;     //500pi/512
   m_sin[501]  =  6'b110110;     //501pi/512
   m_cos[501]  =  6'b110100;     //501pi/512
   m_sin[502]  =  6'b110110;     //502pi/512
   m_cos[502]  =  6'b110100;     //502pi/512
   m_sin[503]  =  6'b110110;     //503pi/512
   m_cos[503]  =  6'b110011;     //503pi/512
   m_sin[504]  =  6'b110110;     //504pi/512
   m_cos[504]  =  6'b110011;     //504pi/512
   m_sin[505]  =  6'b110110;     //505pi/512
   m_cos[505]  =  6'b110011;     //505pi/512
   m_sin[506]  =  6'b110110;     //506pi/512
   m_cos[506]  =  6'b110011;     //506pi/512
   m_sin[507]  =  6'b110110;     //507pi/512
   m_cos[507]  =  6'b110011;     //507pi/512
   m_sin[508]  =  6'b110110;     //508pi/512
   m_cos[508]  =  6'b110011;     //508pi/512
   m_sin[509]  =  6'b110110;     //509pi/512
   m_cos[509]  =  6'b110011;     //509pi/512
   m_sin[510]  =  6'b110110;     //510pi/512
   m_cos[510]  =  6'b110011;     //510pi/512
   m_sin[511]  =  6'b110111;     //511pi/512
   m_cos[511]  =  6'b110011;     //511pi/512
end
endmodule