module  tw_factor_for_9th #(parameter stage_FFT = 2, SIZE =10, word_length_tw = 14) (
    input            clk,
    input            en_rd, 
    input   [stage_FFT-2:0]   rd_ptr_angle,

    output reg  signed [word_length_tw-1:0]   cos_data,
    output reg  signed [word_length_tw-1:0]   sin_data
 );

reg signed [word_length_tw-1:0]  cos  [255:0];
reg signed [word_length_tw-1:0]  sin  [255:0];


//--------------------------------handle read tw factor------------------------------
     always @(posedge clk) begin 
             if (en_rd  ) begin
                  cos_data           <= cos   [rd_ptr_angle];
                  sin_data           <= sin   [rd_ptr_angle];
             end 
        end

//--------------------------------handle read tw factor------------------------------

initial begin
   sin[0]  =  14'b00000000000000;     //0pi/1024
   cos[0]  =  14'b01000000000000;     //0pi/1024
   sin[1]  =  14'b11111111001110;     //4pi/1024
   cos[1]  =  14'b00111111111111;     //4pi/1024
   sin[2]  =  14'b11111110011011;     //8pi/1024
   cos[2]  =  14'b00111111111110;     //8pi/1024
   sin[3]  =  14'b11111101101001;     //12pi/1024
   cos[3]  =  14'b00111111111101;     //12pi/1024
   sin[4]  =  14'b11111100110111;     //16pi/1024
   cos[4]  =  14'b00111111111011;     //16pi/1024
   sin[5]  =  14'b11111100000101;     //20pi/1024
   cos[5]  =  14'b00111111111000;     //20pi/1024
   sin[6]  =  14'b11111011010011;     //24pi/1024
   cos[6]  =  14'b00111111110100;     //24pi/1024
   sin[7]  =  14'b11111010100001;     //28pi/1024
   cos[7]  =  14'b00111111110000;     //28pi/1024
   sin[8]  =  14'b11111001101111;     //32pi/1024
   cos[8]  =  14'b00111111101100;     //32pi/1024
   sin[9]  =  14'b11111000111101;     //36pi/1024
   cos[9]  =  14'b00111111100111;     //36pi/1024
   sin[10]  =  14'b11111000001011;     //40pi/1024
   cos[10]  =  14'b00111111100001;     //40pi/1024
   sin[11]  =  14'b11110111011001;     //44pi/1024
   cos[11]  =  14'b00111111011010;     //44pi/1024
   sin[12]  =  14'b11110110100111;     //48pi/1024
   cos[12]  =  14'b00111111010011;     //48pi/1024
   sin[13]  =  14'b11110101110101;     //52pi/1024
   cos[13]  =  14'b00111111001011;     //52pi/1024
   sin[14]  =  14'b11110101000100;     //56pi/1024
   cos[14]  =  14'b00111111000011;     //56pi/1024
   sin[15]  =  14'b11110100010010;     //60pi/1024
   cos[15]  =  14'b00111110111010;     //60pi/1024
   sin[16]  =  14'b11110011100001;     //64pi/1024
   cos[16]  =  14'b00111110110001;     //64pi/1024
   sin[17]  =  14'b11110010110000;     //68pi/1024
   cos[17]  =  14'b00111110100111;     //68pi/1024
   sin[18]  =  14'b11110001111111;     //72pi/1024
   cos[18]  =  14'b00111110011100;     //72pi/1024
   sin[19]  =  14'b11110001001110;     //76pi/1024
   cos[19]  =  14'b00111110010001;     //76pi/1024
   sin[20]  =  14'b11110000011101;     //80pi/1024
   cos[20]  =  14'b00111110000101;     //80pi/1024
   sin[21]  =  14'b11101111101100;     //84pi/1024
   cos[21]  =  14'b00111101111000;     //84pi/1024
   sin[22]  =  14'b11101110111100;     //88pi/1024
   cos[22]  =  14'b00111101101011;     //88pi/1024
   sin[23]  =  14'b11101110001011;     //92pi/1024
   cos[23]  =  14'b00111101011101;     //92pi/1024
   sin[24]  =  14'b11101101011011;     //96pi/1024
   cos[24]  =  14'b00111101001111;     //96pi/1024
   sin[25]  =  14'b11101100101011;     //100pi/1024
   cos[25]  =  14'b00111101000000;     //100pi/1024
   sin[26]  =  14'b11101011111011;     //104pi/1024
   cos[26]  =  14'b00111100110001;     //104pi/1024
   sin[27]  =  14'b11101011001100;     //108pi/1024
   cos[27]  =  14'b00111100100001;     //108pi/1024
   sin[28]  =  14'b11101010011100;     //112pi/1024
   cos[28]  =  14'b00111100010000;     //112pi/1024
   sin[29]  =  14'b11101001101101;     //116pi/1024
   cos[29]  =  14'b00111011111111;     //116pi/1024
   sin[30]  =  14'b11101000111110;     //120pi/1024
   cos[30]  =  14'b00111011101101;     //120pi/1024
   sin[31]  =  14'b11101000001111;     //124pi/1024
   cos[31]  =  14'b00111011011011;     //124pi/1024
   sin[32]  =  14'b11100111100001;     //128pi/1024
   cos[32]  =  14'b00111011001000;     //128pi/1024
   sin[33]  =  14'b11100110110010;     //132pi/1024
   cos[33]  =  14'b00111010110100;     //132pi/1024
   sin[34]  =  14'b11100110000100;     //136pi/1024
   cos[34]  =  14'b00111010100000;     //136pi/1024
   sin[35]  =  14'b11100101010110;     //140pi/1024
   cos[35]  =  14'b00111010001011;     //140pi/1024
   sin[36]  =  14'b11100100101001;     //144pi/1024
   cos[36]  =  14'b00111001110110;     //144pi/1024
   sin[37]  =  14'b11100011111011;     //148pi/1024
   cos[37]  =  14'b00111001100000;     //148pi/1024
   sin[38]  =  14'b11100011001110;     //152pi/1024
   cos[38]  =  14'b00111001001010;     //152pi/1024
   sin[39]  =  14'b11100010100010;     //156pi/1024
   cos[39]  =  14'b00111000110011;     //156pi/1024
   sin[40]  =  14'b11100001110101;     //160pi/1024
   cos[40]  =  14'b00111000011100;     //160pi/1024
   sin[41]  =  14'b11100001001001;     //164pi/1024
   cos[41]  =  14'b00111000000100;     //164pi/1024
   sin[42]  =  14'b11100000011101;     //168pi/1024
   cos[42]  =  14'b00110111101011;     //168pi/1024
   sin[43]  =  14'b11011111110010;     //172pi/1024
   cos[43]  =  14'b00110111010010;     //172pi/1024
   sin[44]  =  14'b11011111000110;     //176pi/1024
   cos[44]  =  14'b00110110111001;     //176pi/1024
   sin[45]  =  14'b11011110011011;     //180pi/1024
   cos[45]  =  14'b00110110011111;     //180pi/1024
   sin[46]  =  14'b11011101110001;     //184pi/1024
   cos[46]  =  14'b00110110000100;     //184pi/1024
   sin[47]  =  14'b11011101000110;     //188pi/1024
   cos[47]  =  14'b00110101101001;     //188pi/1024
   sin[48]  =  14'b11011100011100;     //192pi/1024
   cos[48]  =  14'b00110101001101;     //192pi/1024
   sin[49]  =  14'b11011011110011;     //196pi/1024
   cos[49]  =  14'b00110100110001;     //196pi/1024
   sin[50]  =  14'b11011011001001;     //200pi/1024
   cos[50]  =  14'b00110100010100;     //200pi/1024
   sin[51]  =  14'b11011010100001;     //204pi/1024
   cos[51]  =  14'b00110011110111;     //204pi/1024
   sin[52]  =  14'b11011001111000;     //208pi/1024
   cos[52]  =  14'b00110011011001;     //208pi/1024
   sin[53]  =  14'b11011001010000;     //212pi/1024
   cos[53]  =  14'b00110010111011;     //212pi/1024
   sin[54]  =  14'b11011000101000;     //216pi/1024
   cos[54]  =  14'b00110010011101;     //216pi/1024
   sin[55]  =  14'b11011000000001;     //220pi/1024
   cos[55]  =  14'b00110001111101;     //220pi/1024
   sin[56]  =  14'b11010111011010;     //224pi/1024
   cos[56]  =  14'b00110001011110;     //224pi/1024
   sin[57]  =  14'b11010110110011;     //228pi/1024
   cos[57]  =  14'b00110000111110;     //228pi/1024
   sin[58]  =  14'b11010110001101;     //232pi/1024
   cos[58]  =  14'b00110000011101;     //232pi/1024
   sin[59]  =  14'b11010101100111;     //236pi/1024
   cos[59]  =  14'b00101111111100;     //236pi/1024
   sin[60]  =  14'b11010101000001;     //240pi/1024
   cos[60]  =  14'b00101111011010;     //240pi/1024
   sin[61]  =  14'b11010100011100;     //244pi/1024
   cos[61]  =  14'b00101110111000;     //244pi/1024
   sin[62]  =  14'b11010011111000;     //248pi/1024
   cos[62]  =  14'b00101110010110;     //248pi/1024
   sin[63]  =  14'b11010011010011;     //252pi/1024
   cos[63]  =  14'b00101101110011;     //252pi/1024
   sin[64]  =  14'b11010010110000;     //256pi/1024
   cos[64]  =  14'b00101101010000;     //256pi/1024
   sin[65]  =  14'b11010010001100;     //260pi/1024
   cos[65]  =  14'b00101100101100;     //260pi/1024
   sin[66]  =  14'b11010001101001;     //264pi/1024
   cos[66]  =  14'b00101100001000;     //264pi/1024
   sin[67]  =  14'b11010001000111;     //268pi/1024
   cos[67]  =  14'b00101011100011;     //268pi/1024
   sin[68]  =  14'b11010000100101;     //272pi/1024
   cos[68]  =  14'b00101010111110;     //272pi/1024
   sin[69]  =  14'b11010000000100;     //276pi/1024
   cos[69]  =  14'b00101010011001;     //276pi/1024
   sin[70]  =  14'b11001111100010;     //280pi/1024
   cos[70]  =  14'b00101001110011;     //280pi/1024
   sin[71]  =  14'b11001111000010;     //284pi/1024
   cos[71]  =  14'b00101001001101;     //284pi/1024
   sin[72]  =  14'b11001110100010;     //288pi/1024
   cos[72]  =  14'b00101000100110;     //288pi/1024
   sin[73]  =  14'b11001110000010;     //292pi/1024
   cos[73]  =  14'b00100111111111;     //292pi/1024
   sin[74]  =  14'b11001101100011;     //296pi/1024
   cos[74]  =  14'b00100111010111;     //296pi/1024
   sin[75]  =  14'b11001101000100;     //300pi/1024
   cos[75]  =  14'b00100110110000;     //300pi/1024
   sin[76]  =  14'b11001100100110;     //304pi/1024
   cos[76]  =  14'b00100110000111;     //304pi/1024
   sin[77]  =  14'b11001100001000;     //308pi/1024
   cos[77]  =  14'b00100101011111;     //308pi/1024
   sin[78]  =  14'b11001011101011;     //312pi/1024
   cos[78]  =  14'b00100100110110;     //312pi/1024
   sin[79]  =  14'b11001011001110;     //316pi/1024
   cos[79]  =  14'b00100100001101;     //316pi/1024
   sin[80]  =  14'b11001010110010;     //320pi/1024
   cos[80]  =  14'b00100011100011;     //320pi/1024
   sin[81]  =  14'b11001010010111;     //324pi/1024
   cos[81]  =  14'b00100010111001;     //324pi/1024
   sin[82]  =  14'b11001001111011;     //328pi/1024
   cos[82]  =  14'b00100010001111;     //328pi/1024
   sin[83]  =  14'b11001001100001;     //332pi/1024
   cos[83]  =  14'b00100001100100;     //332pi/1024
   sin[84]  =  14'b11001001000111;     //336pi/1024
   cos[84]  =  14'b00100000111001;     //336pi/1024
   sin[85]  =  14'b11001000101101;     //340pi/1024
   cos[85]  =  14'b00100000001110;     //340pi/1024
   sin[86]  =  14'b11001000010100;     //344pi/1024
   cos[86]  =  14'b00011111100010;     //344pi/1024
   sin[87]  =  14'b11000111111100;     //348pi/1024
   cos[87]  =  14'b00011110110111;     //348pi/1024
   sin[88]  =  14'b11000111100100;     //352pi/1024
   cos[88]  =  14'b00011110001010;     //352pi/1024
   sin[89]  =  14'b11000111001100;     //356pi/1024
   cos[89]  =  14'b00011101011110;     //356pi/1024
   sin[90]  =  14'b11000110110101;     //360pi/1024
   cos[90]  =  14'b00011100110001;     //360pi/1024
   sin[91]  =  14'b11000110011111;     //364pi/1024
   cos[91]  =  14'b00011100000100;     //364pi/1024
   sin[92]  =  14'b11000110001001;     //368pi/1024
   cos[92]  =  14'b00011011010111;     //368pi/1024
   sin[93]  =  14'b11000101110100;     //372pi/1024
   cos[93]  =  14'b00011010101001;     //372pi/1024
   sin[94]  =  14'b11000101011111;     //376pi/1024
   cos[94]  =  14'b00011001111011;     //376pi/1024
   sin[95]  =  14'b11000101001011;     //380pi/1024
   cos[95]  =  14'b00011001001101;     //380pi/1024
   sin[96]  =  14'b11000100111000;     //384pi/1024
   cos[96]  =  14'b00011000011111;     //384pi/1024
   sin[97]  =  14'b11000100100101;     //388pi/1024
   cos[97]  =  14'b00010111110000;     //388pi/1024
   sin[98]  =  14'b11000100010010;     //392pi/1024
   cos[98]  =  14'b00010111000010;     //392pi/1024
   sin[99]  =  14'b11000100000001;     //396pi/1024
   cos[99]  =  14'b00010110010011;     //396pi/1024
   sin[100]  =  14'b11000011101111;     //400pi/1024
   cos[100]  =  14'b00010101100011;     //400pi/1024
   sin[101]  =  14'b11000011011111;     //404pi/1024
   cos[101]  =  14'b00010100110100;     //404pi/1024
   sin[102]  =  14'b11000011001111;     //408pi/1024
   cos[102]  =  14'b00010100000100;     //408pi/1024
   sin[103]  =  14'b11000010111111;     //412pi/1024
   cos[103]  =  14'b00010011010101;     //412pi/1024
   sin[104]  =  14'b11000010110000;     //416pi/1024
   cos[104]  =  14'b00010010100101;     //416pi/1024
   sin[105]  =  14'b11000010100010;     //420pi/1024
   cos[105]  =  14'b00010001110100;     //420pi/1024
   sin[106]  =  14'b11000010010100;     //424pi/1024
   cos[106]  =  14'b00010001000100;     //424pi/1024
   sin[107]  =  14'b11000010000111;     //428pi/1024
   cos[107]  =  14'b00010000010011;     //428pi/1024
   sin[108]  =  14'b11000001111011;     //432pi/1024
   cos[108]  =  14'b00001111100011;     //432pi/1024
   sin[109]  =  14'b11000001101111;     //436pi/1024
   cos[109]  =  14'b00001110110010;     //436pi/1024
   sin[110]  =  14'b11000001100100;     //440pi/1024
   cos[110]  =  14'b00001110000001;     //440pi/1024
   sin[111]  =  14'b11000001011001;     //444pi/1024
   cos[111]  =  14'b00001101010000;     //444pi/1024
   sin[112]  =  14'b11000001001111;     //448pi/1024
   cos[112]  =  14'b00001100011111;     //448pi/1024
   sin[113]  =  14'b11000001000101;     //452pi/1024
   cos[113]  =  14'b00001011101101;     //452pi/1024
   sin[114]  =  14'b11000000111100;     //456pi/1024
   cos[114]  =  14'b00001010111100;     //456pi/1024
   sin[115]  =  14'b11000000110100;     //460pi/1024
   cos[115]  =  14'b00001010001010;     //460pi/1024
   sin[116]  =  14'b11000000101100;     //464pi/1024
   cos[116]  =  14'b00001001011001;     //464pi/1024
   sin[117]  =  14'b11000000100101;     //468pi/1024
   cos[117]  =  14'b00001000100111;     //468pi/1024
   sin[118]  =  14'b11000000011111;     //472pi/1024
   cos[118]  =  14'b00000111110101;     //472pi/1024
   sin[119]  =  14'b11000000011001;     //476pi/1024
   cos[119]  =  14'b00000111000011;     //476pi/1024
   sin[120]  =  14'b11000000010100;     //480pi/1024
   cos[120]  =  14'b00000110010001;     //480pi/1024
   sin[121]  =  14'b11000000001111;     //484pi/1024
   cos[121]  =  14'b00000101011111;     //484pi/1024
   sin[122]  =  14'b11000000001011;     //488pi/1024
   cos[122]  =  14'b00000100101101;     //488pi/1024
   sin[123]  =  14'b11000000001000;     //492pi/1024
   cos[123]  =  14'b00000011111011;     //492pi/1024
   sin[124]  =  14'b11000000000101;     //496pi/1024
   cos[124]  =  14'b00000011001000;     //496pi/1024
   sin[125]  =  14'b11000000000011;     //500pi/1024
   cos[125]  =  14'b00000010010110;     //500pi/1024
   sin[126]  =  14'b11000000000001;     //504pi/1024
   cos[126]  =  14'b00000001100100;     //504pi/1024
   sin[127]  =  14'b11000000000000;     //508pi/1024
   cos[127]  =  14'b00000000110010;     //508pi/1024
   sin[128]  =  14'b11000000000000;     //512pi/1024
   cos[128]  =  14'b00000000000000;     //512pi/1024
   sin[129]  =  14'b11000000000000;     //516pi/1024
   cos[129]  =  14'b11111111001110;     //516pi/1024
   sin[130]  =  14'b11000000000001;     //520pi/1024
   cos[130]  =  14'b11111110011011;     //520pi/1024
   sin[131]  =  14'b11000000000011;     //524pi/1024
   cos[131]  =  14'b11111101101001;     //524pi/1024
   sin[132]  =  14'b11000000000101;     //528pi/1024
   cos[132]  =  14'b11111100110111;     //528pi/1024
   sin[133]  =  14'b11000000001000;     //532pi/1024
   cos[133]  =  14'b11111100000101;     //532pi/1024
   sin[134]  =  14'b11000000001011;     //536pi/1024
   cos[134]  =  14'b11111011010011;     //536pi/1024
   sin[135]  =  14'b11000000001111;     //540pi/1024
   cos[135]  =  14'b11111010100001;     //540pi/1024
   sin[136]  =  14'b11000000010100;     //544pi/1024
   cos[136]  =  14'b11111001101111;     //544pi/1024
   sin[137]  =  14'b11000000011001;     //548pi/1024
   cos[137]  =  14'b11111000111101;     //548pi/1024
   sin[138]  =  14'b11000000011111;     //552pi/1024
   cos[138]  =  14'b11111000001011;     //552pi/1024
   sin[139]  =  14'b11000000100101;     //556pi/1024
   cos[139]  =  14'b11110111011001;     //556pi/1024
   sin[140]  =  14'b11000000101100;     //560pi/1024
   cos[140]  =  14'b11110110100111;     //560pi/1024
   sin[141]  =  14'b11000000110100;     //564pi/1024
   cos[141]  =  14'b11110101110101;     //564pi/1024
   sin[142]  =  14'b11000000111100;     //568pi/1024
   cos[142]  =  14'b11110101000100;     //568pi/1024
   sin[143]  =  14'b11000001000101;     //572pi/1024
   cos[143]  =  14'b11110100010010;     //572pi/1024
   sin[144]  =  14'b11000001001111;     //576pi/1024
   cos[144]  =  14'b11110011100001;     //576pi/1024
   sin[145]  =  14'b11000001011001;     //580pi/1024
   cos[145]  =  14'b11110010110000;     //580pi/1024
   sin[146]  =  14'b11000001100100;     //584pi/1024
   cos[146]  =  14'b11110001111111;     //584pi/1024
   sin[147]  =  14'b11000001101111;     //588pi/1024
   cos[147]  =  14'b11110001001110;     //588pi/1024
   sin[148]  =  14'b11000001111011;     //592pi/1024
   cos[148]  =  14'b11110000011101;     //592pi/1024
   sin[149]  =  14'b11000010000111;     //596pi/1024
   cos[149]  =  14'b11101111101100;     //596pi/1024
   sin[150]  =  14'b11000010010100;     //600pi/1024
   cos[150]  =  14'b11101110111100;     //600pi/1024
   sin[151]  =  14'b11000010100010;     //604pi/1024
   cos[151]  =  14'b11101110001011;     //604pi/1024
   sin[152]  =  14'b11000010110000;     //608pi/1024
   cos[152]  =  14'b11101101011011;     //608pi/1024
   sin[153]  =  14'b11000010111111;     //612pi/1024
   cos[153]  =  14'b11101100101011;     //612pi/1024
   sin[154]  =  14'b11000011001111;     //616pi/1024
   cos[154]  =  14'b11101011111011;     //616pi/1024
   sin[155]  =  14'b11000011011111;     //620pi/1024
   cos[155]  =  14'b11101011001100;     //620pi/1024
   sin[156]  =  14'b11000011101111;     //624pi/1024
   cos[156]  =  14'b11101010011100;     //624pi/1024
   sin[157]  =  14'b11000100000001;     //628pi/1024
   cos[157]  =  14'b11101001101101;     //628pi/1024
   sin[158]  =  14'b11000100010010;     //632pi/1024
   cos[158]  =  14'b11101000111110;     //632pi/1024
   sin[159]  =  14'b11000100100101;     //636pi/1024
   cos[159]  =  14'b11101000001111;     //636pi/1024
   sin[160]  =  14'b11000100111000;     //640pi/1024
   cos[160]  =  14'b11100111100001;     //640pi/1024
   sin[161]  =  14'b11000101001011;     //644pi/1024
   cos[161]  =  14'b11100110110010;     //644pi/1024
   sin[162]  =  14'b11000101011111;     //648pi/1024
   cos[162]  =  14'b11100110000100;     //648pi/1024
   sin[163]  =  14'b11000101110100;     //652pi/1024
   cos[163]  =  14'b11100101010110;     //652pi/1024
   sin[164]  =  14'b11000110001001;     //656pi/1024
   cos[164]  =  14'b11100100101001;     //656pi/1024
   sin[165]  =  14'b11000110011111;     //660pi/1024
   cos[165]  =  14'b11100011111011;     //660pi/1024
   sin[166]  =  14'b11000110110101;     //664pi/1024
   cos[166]  =  14'b11100011001110;     //664pi/1024
   sin[167]  =  14'b11000111001100;     //668pi/1024
   cos[167]  =  14'b11100010100010;     //668pi/1024
   sin[168]  =  14'b11000111100100;     //672pi/1024
   cos[168]  =  14'b11100001110101;     //672pi/1024
   sin[169]  =  14'b11000111111100;     //676pi/1024
   cos[169]  =  14'b11100001001001;     //676pi/1024
   sin[170]  =  14'b11001000010100;     //680pi/1024
   cos[170]  =  14'b11100000011101;     //680pi/1024
   sin[171]  =  14'b11001000101101;     //684pi/1024
   cos[171]  =  14'b11011111110010;     //684pi/1024
   sin[172]  =  14'b11001001000111;     //688pi/1024
   cos[172]  =  14'b11011111000110;     //688pi/1024
   sin[173]  =  14'b11001001100001;     //692pi/1024
   cos[173]  =  14'b11011110011011;     //692pi/1024
   sin[174]  =  14'b11001001111011;     //696pi/1024
   cos[174]  =  14'b11011101110001;     //696pi/1024
   sin[175]  =  14'b11001010010111;     //700pi/1024
   cos[175]  =  14'b11011101000110;     //700pi/1024
   sin[176]  =  14'b11001010110010;     //704pi/1024
   cos[176]  =  14'b11011100011100;     //704pi/1024
   sin[177]  =  14'b11001011001110;     //708pi/1024
   cos[177]  =  14'b11011011110011;     //708pi/1024
   sin[178]  =  14'b11001011101011;     //712pi/1024
   cos[178]  =  14'b11011011001001;     //712pi/1024
   sin[179]  =  14'b11001100001000;     //716pi/1024
   cos[179]  =  14'b11011010100001;     //716pi/1024
   sin[180]  =  14'b11001100100110;     //720pi/1024
   cos[180]  =  14'b11011001111000;     //720pi/1024
   sin[181]  =  14'b11001101000100;     //724pi/1024
   cos[181]  =  14'b11011001010000;     //724pi/1024
   sin[182]  =  14'b11001101100011;     //728pi/1024
   cos[182]  =  14'b11011000101000;     //728pi/1024
   sin[183]  =  14'b11001110000010;     //732pi/1024
   cos[183]  =  14'b11011000000001;     //732pi/1024
   sin[184]  =  14'b11001110100010;     //736pi/1024
   cos[184]  =  14'b11010111011010;     //736pi/1024
   sin[185]  =  14'b11001111000010;     //740pi/1024
   cos[185]  =  14'b11010110110011;     //740pi/1024
   sin[186]  =  14'b11001111100010;     //744pi/1024
   cos[186]  =  14'b11010110001101;     //744pi/1024
   sin[187]  =  14'b11010000000100;     //748pi/1024
   cos[187]  =  14'b11010101100111;     //748pi/1024
   sin[188]  =  14'b11010000100101;     //752pi/1024
   cos[188]  =  14'b11010101000001;     //752pi/1024
   sin[189]  =  14'b11010001000111;     //756pi/1024
   cos[189]  =  14'b11010100011100;     //756pi/1024
   sin[190]  =  14'b11010001101001;     //760pi/1024
   cos[190]  =  14'b11010011111000;     //760pi/1024
   sin[191]  =  14'b11010010001100;     //764pi/1024
   cos[191]  =  14'b11010011010011;     //764pi/1024
   sin[192]  =  14'b11010010110000;     //768pi/1024
   cos[192]  =  14'b11010010110000;     //768pi/1024
   sin[193]  =  14'b11010011010011;     //772pi/1024
   cos[193]  =  14'b11010010001100;     //772pi/1024
   sin[194]  =  14'b11010011111000;     //776pi/1024
   cos[194]  =  14'b11010001101001;     //776pi/1024
   sin[195]  =  14'b11010100011100;     //780pi/1024
   cos[195]  =  14'b11010001000111;     //780pi/1024
   sin[196]  =  14'b11010101000001;     //784pi/1024
   cos[196]  =  14'b11010000100101;     //784pi/1024
   sin[197]  =  14'b11010101100111;     //788pi/1024
   cos[197]  =  14'b11010000000100;     //788pi/1024
   sin[198]  =  14'b11010110001101;     //792pi/1024
   cos[198]  =  14'b11001111100010;     //792pi/1024
   sin[199]  =  14'b11010110110011;     //796pi/1024
   cos[199]  =  14'b11001111000010;     //796pi/1024
   sin[200]  =  14'b11010111011010;     //800pi/1024
   cos[200]  =  14'b11001110100010;     //800pi/1024
   sin[201]  =  14'b11011000000001;     //804pi/1024
   cos[201]  =  14'b11001110000010;     //804pi/1024
   sin[202]  =  14'b11011000101000;     //808pi/1024
   cos[202]  =  14'b11001101100011;     //808pi/1024
   sin[203]  =  14'b11011001010000;     //812pi/1024
   cos[203]  =  14'b11001101000100;     //812pi/1024
   sin[204]  =  14'b11011001111000;     //816pi/1024
   cos[204]  =  14'b11001100100110;     //816pi/1024
   sin[205]  =  14'b11011010100001;     //820pi/1024
   cos[205]  =  14'b11001100001000;     //820pi/1024
   sin[206]  =  14'b11011011001001;     //824pi/1024
   cos[206]  =  14'b11001011101011;     //824pi/1024
   sin[207]  =  14'b11011011110011;     //828pi/1024
   cos[207]  =  14'b11001011001110;     //828pi/1024
   sin[208]  =  14'b11011100011100;     //832pi/1024
   cos[208]  =  14'b11001010110010;     //832pi/1024
   sin[209]  =  14'b11011101000110;     //836pi/1024
   cos[209]  =  14'b11001010010111;     //836pi/1024
   sin[210]  =  14'b11011101110001;     //840pi/1024
   cos[210]  =  14'b11001001111011;     //840pi/1024
   sin[211]  =  14'b11011110011011;     //844pi/1024
   cos[211]  =  14'b11001001100001;     //844pi/1024
   sin[212]  =  14'b11011111000110;     //848pi/1024
   cos[212]  =  14'b11001001000111;     //848pi/1024
   sin[213]  =  14'b11011111110010;     //852pi/1024
   cos[213]  =  14'b11001000101101;     //852pi/1024
   sin[214]  =  14'b11100000011101;     //856pi/1024
   cos[214]  =  14'b11001000010100;     //856pi/1024
   sin[215]  =  14'b11100001001001;     //860pi/1024
   cos[215]  =  14'b11000111111100;     //860pi/1024
   sin[216]  =  14'b11100001110101;     //864pi/1024
   cos[216]  =  14'b11000111100100;     //864pi/1024
   sin[217]  =  14'b11100010100010;     //868pi/1024
   cos[217]  =  14'b11000111001100;     //868pi/1024
   sin[218]  =  14'b11100011001110;     //872pi/1024
   cos[218]  =  14'b11000110110101;     //872pi/1024
   sin[219]  =  14'b11100011111011;     //876pi/1024
   cos[219]  =  14'b11000110011111;     //876pi/1024
   sin[220]  =  14'b11100100101001;     //880pi/1024
   cos[220]  =  14'b11000110001001;     //880pi/1024
   sin[221]  =  14'b11100101010110;     //884pi/1024
   cos[221]  =  14'b11000101110100;     //884pi/1024
   sin[222]  =  14'b11100110000100;     //888pi/1024
   cos[222]  =  14'b11000101011111;     //888pi/1024
   sin[223]  =  14'b11100110110010;     //892pi/1024
   cos[223]  =  14'b11000101001011;     //892pi/1024
   sin[224]  =  14'b11100111100001;     //896pi/1024
   cos[224]  =  14'b11000100111000;     //896pi/1024
   sin[225]  =  14'b11101000001111;     //900pi/1024
   cos[225]  =  14'b11000100100101;     //900pi/1024
   sin[226]  =  14'b11101000111110;     //904pi/1024
   cos[226]  =  14'b11000100010010;     //904pi/1024
   sin[227]  =  14'b11101001101101;     //908pi/1024
   cos[227]  =  14'b11000100000001;     //908pi/1024
   sin[228]  =  14'b11101010011100;     //912pi/1024
   cos[228]  =  14'b11000011101111;     //912pi/1024
   sin[229]  =  14'b11101011001100;     //916pi/1024
   cos[229]  =  14'b11000011011111;     //916pi/1024
   sin[230]  =  14'b11101011111011;     //920pi/1024
   cos[230]  =  14'b11000011001111;     //920pi/1024
   sin[231]  =  14'b11101100101011;     //924pi/1024
   cos[231]  =  14'b11000010111111;     //924pi/1024
   sin[232]  =  14'b11101101011011;     //928pi/1024
   cos[232]  =  14'b11000010110000;     //928pi/1024
   sin[233]  =  14'b11101110001011;     //932pi/1024
   cos[233]  =  14'b11000010100010;     //932pi/1024
   sin[234]  =  14'b11101110111100;     //936pi/1024
   cos[234]  =  14'b11000010010100;     //936pi/1024
   sin[235]  =  14'b11101111101100;     //940pi/1024
   cos[235]  =  14'b11000010000111;     //940pi/1024
   sin[236]  =  14'b11110000011101;     //944pi/1024
   cos[236]  =  14'b11000001111011;     //944pi/1024
   sin[237]  =  14'b11110001001110;     //948pi/1024
   cos[237]  =  14'b11000001101111;     //948pi/1024
   sin[238]  =  14'b11110001111111;     //952pi/1024
   cos[238]  =  14'b11000001100100;     //952pi/1024
   sin[239]  =  14'b11110010110000;     //956pi/1024
   cos[239]  =  14'b11000001011001;     //956pi/1024
   sin[240]  =  14'b11110011100001;     //960pi/1024
   cos[240]  =  14'b11000001001111;     //960pi/1024
   sin[241]  =  14'b11110100010010;     //964pi/1024
   cos[241]  =  14'b11000001000101;     //964pi/1024
   sin[242]  =  14'b11110101000100;     //968pi/1024
   cos[242]  =  14'b11000000111100;     //968pi/1024
   sin[243]  =  14'b11110101110101;     //972pi/1024
   cos[243]  =  14'b11000000110100;     //972pi/1024
   sin[244]  =  14'b11110110100111;     //976pi/1024
   cos[244]  =  14'b11000000101100;     //976pi/1024
   sin[245]  =  14'b11110111011001;     //980pi/1024
   cos[245]  =  14'b11000000100101;     //980pi/1024
   sin[246]  =  14'b11111000001011;     //984pi/1024
   cos[246]  =  14'b11000000011111;     //984pi/1024
   sin[247]  =  14'b11111000111101;     //988pi/1024
   cos[247]  =  14'b11000000011001;     //988pi/1024
   sin[248]  =  14'b11111001101111;     //992pi/1024
   cos[248]  =  14'b11000000010100;     //992pi/1024
   sin[249]  =  14'b11111010100001;     //996pi/1024
   cos[249]  =  14'b11000000001111;     //996pi/1024
   sin[250]  =  14'b11111011010011;     //1000pi/1024
   cos[250]  =  14'b11000000001011;     //1000pi/1024
   sin[251]  =  14'b11111100000101;     //1004pi/1024
   cos[251]  =  14'b11000000001000;     //1004pi/1024
   sin[252]  =  14'b11111100110111;     //1008pi/1024
   cos[252]  =  14'b11000000000101;     //1008pi/1024
   sin[253]  =  14'b11111101101001;     //1012pi/1024
   cos[253]  =  14'b11000000000011;     //1012pi/1024
   sin[254]  =  14'b11111110011011;     //1016pi/1024
   cos[254]  =  14'b11000000000001;     //1016pi/1024
   sin[255]  =  14'b11111111001110;     //1020pi/1024
   cos[255]  =  14'b11000000000000;     //1020pi/1024
end
endmodule